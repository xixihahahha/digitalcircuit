`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2023/11/09 15:05:05
// Design Name: 
// Module Name: key_Create
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module SM4(
    input [127:0] MK,
    input [127:0] plain,
    output reg [127:0] cipher
    );
    
    reg [31:0] FK [0:3];
    reg [31:0] CK [0:31];
    
    reg [31:0] RK [0:35];
    reg [31:0] text [0:35];
    reg [31:0] num = 0;
    initial begin
        FK[0] = 0'ha3b1bac6;
        FK[1] = 0'h56aa3350;
        FK[2] = 0'h677d9197;
        FK[3] = 0'hb27022dc;
        
        CK[0] = 0'h00070e15;
        CK[1] = 0'h1c232a31;
        CK[2] = 0'h383f464d;
        CK[3] = 0'h545b6269;
        CK[4] = 0'h70777e85;
        CK[5] = 0'h8c939aa1;
        CK[6] = 0'ha8afb6bd;
        CK[7] = 0'hc4cbd2d9;
        CK[8] = 0'he0e7eef5;
        CK[9] = 0'hfc030a11;
        CK[10] = 0'h181f262d;
        CK[11] = 0'h343b4249;
        CK[12] = 0'h50575e65;
        CK[13] = 0'h6c737a81;
        CK[14] = 0'h888f969d;
        CK[15] = 0'ha4abb2b9;
        CK[16] = 0'hc0c7ced5;
        CK[17] = 0'hdce3eaf1;
        CK[18] = 0'hf8ff060d;
        CK[19] = 0'h141b2229;
        CK[20] = 0'h30373e45;
        CK[21] = 0'h4c535a61;
        CK[22] = 0'h686f767d;
        CK[23] = 0'h848b9299;
        CK[24] = 0'ha0a7aeb5;
        CK[25] = 0'hbcc3cad1;
        CK[26] = 0'hd8dfe6ed;
        CK[27] = 0'hf4fb0209;
        CK[28] = 0'h10171e25;
        CK[29] = 0'h2c333a41;
        CK[30] = 0'h484f565d;
        CK[31] = 0'h646b7279;
    end
    
    integer i;
    always @(*) begin
    RK[0] = MK[127:96] ^ FK[0];
    RK[1] = MK[95:64] ^ FK[1];
    RK[2] = MK[63:32] ^ FK[2];
    RK[3] = MK[31:0] ^ FK[3];
    for(i = 0; i < 32; i = i + 1) begin
        num = RK[i+1] ^ RK[i+2] ^ RK[i+3] ^ CK[i];
        
        case(num[7:0])
	8'h00: num[7:0] = 8'hd6;
	8'h01: num[7:0] = 8'h90;
	8'h02: num[7:0] = 8'he9;
	8'h03: num[7:0] = 8'hfe;
	8'h04: num[7:0] = 8'hcc;
	8'h05: num[7:0] = 8'he1;
	8'h06: num[7:0] = 8'h3d;
	8'h07: num[7:0] = 8'hb7;
	8'h08: num[7:0] = 8'h16;
	8'h09: num[7:0] = 8'hb6;
	8'h0a: num[7:0] = 8'h14;
	8'h0b: num[7:0] = 8'hc2;
	8'h0c: num[7:0] = 8'h28;
	8'h0d: num[7:0] = 8'hfb;
	8'h0e: num[7:0] = 8'h2c;
	8'h0f: num[7:0] = 8'h05;
	8'h10: num[7:0] = 8'h2b;
	8'h11: num[7:0] = 8'h67;
	8'h12: num[7:0] = 8'h9a;
	8'h13: num[7:0] = 8'h76;
	8'h14: num[7:0] = 8'h2a;
	8'h15: num[7:0] = 8'hbe;
	8'h16: num[7:0] = 8'h04;
	8'h17: num[7:0] = 8'hc3;
	8'h18: num[7:0] = 8'haa;
	8'h19: num[7:0] = 8'h44;
	8'h1a: num[7:0] = 8'h13;
	8'h1b: num[7:0] = 8'h26;
	8'h1c: num[7:0] = 8'h49;
	8'h1d: num[7:0] = 8'h86;
	8'h1e: num[7:0] = 8'h06;
	8'h1f: num[7:0] = 8'h99;
	8'h20: num[7:0] = 8'h9c;
	8'h21: num[7:0] = 8'h42;
	8'h22: num[7:0] = 8'h50;
	8'h23: num[7:0] = 8'hf4;
	8'h24: num[7:0] = 8'h91;
	8'h25: num[7:0] = 8'hef;
	8'h26: num[7:0] = 8'h98;
	8'h27: num[7:0] = 8'h7a;
	8'h28: num[7:0] = 8'h33;
	8'h29: num[7:0] = 8'h54;
	8'h2a: num[7:0] = 8'h0b;
	8'h2b: num[7:0] = 8'h43;
	8'h2c: num[7:0] = 8'hed;
	8'h2d: num[7:0] = 8'hcf;
	8'h2e: num[7:0] = 8'hac;
	8'h2f: num[7:0] = 8'h62;
	8'h30: num[7:0] = 8'he4;
	8'h31: num[7:0] = 8'hb3;
	8'h32: num[7:0] = 8'h1c;
	8'h33: num[7:0] = 8'ha9;
	8'h34: num[7:0] = 8'hc9;
	8'h35: num[7:0] = 8'h08;
	8'h36: num[7:0] = 8'he8;
	8'h37: num[7:0] = 8'h95;
	8'h38: num[7:0] = 8'h80;
	8'h39: num[7:0] = 8'hdf;
	8'h3a: num[7:0] = 8'h94;
	8'h3b: num[7:0] = 8'hfa;
	8'h3c: num[7:0] = 8'h75;
	8'h3d: num[7:0] = 8'h8f;
	8'h3e: num[7:0] = 8'h3f;
	8'h3f: num[7:0] = 8'ha6;
	8'h40: num[7:0] = 8'h47;
	8'h41: num[7:0] = 8'h07;
	8'h42: num[7:0] = 8'ha7;
	8'h43: num[7:0] = 8'hfc;
	8'h44: num[7:0] = 8'hf3;
	8'h45: num[7:0] = 8'h73;
	8'h46: num[7:0] = 8'h17;
	8'h47: num[7:0] = 8'hba;
	8'h48: num[7:0] = 8'h83;
	8'h49: num[7:0] = 8'h59;
	8'h4a: num[7:0] = 8'h3c;
	8'h4b: num[7:0] = 8'h19;
	8'h4c: num[7:0] = 8'he6;
	8'h4d: num[7:0] = 8'h85;
	8'h4e: num[7:0] = 8'h4f;
	8'h4f: num[7:0] = 8'ha8;
	8'h50: num[7:0] = 8'h68;
	8'h51: num[7:0] = 8'h6b;
	8'h52: num[7:0] = 8'h81;
	8'h53: num[7:0] = 8'hb2;
	8'h54: num[7:0] = 8'h71;
	8'h55: num[7:0] = 8'h64;
	8'h56: num[7:0] = 8'hda;
	8'h57: num[7:0] = 8'h8b;
	8'h58: num[7:0] = 8'hf8;
	8'h59: num[7:0] = 8'heb;
	8'h5a: num[7:0] = 8'h0f;
	8'h5b: num[7:0] = 8'h4b;
	8'h5c: num[7:0] = 8'h70;
	8'h5d: num[7:0] = 8'h56;
	8'h5e: num[7:0] = 8'h9d;
	8'h5f: num[7:0] = 8'h35;
	8'h60: num[7:0] = 8'h1e;
	8'h61: num[7:0] = 8'h24;
	8'h62: num[7:0] = 8'h0e;
	8'h63: num[7:0] = 8'h5e;
	8'h64: num[7:0] = 8'h63;
	8'h65: num[7:0] = 8'h58;
	8'h66: num[7:0] = 8'hd1;
	8'h67: num[7:0] = 8'ha2;
	8'h68: num[7:0] = 8'h25;
	8'h69: num[7:0] = 8'h22;
	8'h6a: num[7:0] = 8'h7c;
	8'h6b: num[7:0] = 8'h3b;
	8'h6c: num[7:0] = 8'h01;
	8'h6d: num[7:0] = 8'h21;
	8'h6e: num[7:0] = 8'h78;
	8'h6f: num[7:0] = 8'h87;
	8'h70: num[7:0] = 8'hd4;
	8'h71: num[7:0] = 8'h00;
	8'h72: num[7:0] = 8'h46;
	8'h73: num[7:0] = 8'h57;
	8'h74: num[7:0] = 8'h9f;
	8'h75: num[7:0] = 8'hd3;
	8'h76: num[7:0] = 8'h27;
	8'h77: num[7:0] = 8'h52;
	8'h78: num[7:0] = 8'h4c;
	8'h79: num[7:0] = 8'h36;
	8'h7a: num[7:0] = 8'h02;
	8'h7b: num[7:0] = 8'he7;
	8'h7c: num[7:0] = 8'ha0;
	8'h7d: num[7:0] = 8'hc4;
	8'h7e: num[7:0] = 8'hc8;
	8'h7f: num[7:0] = 8'h9e;
	8'h80: num[7:0] = 8'hea;
	8'h81: num[7:0] = 8'hbf;
	8'h82: num[7:0] = 8'h8a;
	8'h83: num[7:0] = 8'hd2;
	8'h84: num[7:0] = 8'h40;
	8'h85: num[7:0] = 8'hc7;
	8'h86: num[7:0] = 8'h38;
	8'h87: num[7:0] = 8'hb5;
	8'h88: num[7:0] = 8'ha3;
	8'h89: num[7:0] = 8'hf7;
	8'h8a: num[7:0] = 8'hf2;
	8'h8b: num[7:0] = 8'hce;
	8'h8c: num[7:0] = 8'hf9;
	8'h8d: num[7:0] = 8'h61;
	8'h8e: num[7:0] = 8'h15;
	8'h8f: num[7:0] = 8'ha1;
	8'h90: num[7:0] = 8'he0;
	8'h91: num[7:0] = 8'hae;
	8'h92: num[7:0] = 8'h5d;
	8'h93: num[7:0] = 8'ha4;
	8'h94: num[7:0] = 8'h9b;
	8'h95: num[7:0] = 8'h34;
	8'h96: num[7:0] = 8'h1a;
	8'h97: num[7:0] = 8'h55;
	8'h98: num[7:0] = 8'had;
	8'h99: num[7:0] = 8'h93;
	8'h9a: num[7:0] = 8'h32;
	8'h9b: num[7:0] = 8'h30;
	8'h9c: num[7:0] = 8'hf5;
	8'h9d: num[7:0] = 8'h8c;
	8'h9e: num[7:0] = 8'hb1;
	8'h9f: num[7:0] = 8'he3;
	8'ha0: num[7:0] = 8'h1d;
	8'ha1: num[7:0] = 8'hf6;
	8'ha2: num[7:0] = 8'he2;
	8'ha3: num[7:0] = 8'h2e;
	8'ha4: num[7:0] = 8'h82;
	8'ha5: num[7:0] = 8'h66;
	8'ha6: num[7:0] = 8'hca;
	8'ha7: num[7:0] = 8'h60;
	8'ha8: num[7:0] = 8'hc0;
	8'ha9: num[7:0] = 8'h29;
	8'haa: num[7:0] = 8'h23;
	8'hab: num[7:0] = 8'hab;
	8'hac: num[7:0] = 8'h0d;
	8'had: num[7:0] = 8'h53;
	8'hae: num[7:0] = 8'h4e;
	8'haf: num[7:0] = 8'h6f;
	8'hb0: num[7:0] = 8'hd5;
	8'hb1: num[7:0] = 8'hdb;
	8'hb2: num[7:0] = 8'h37;
	8'hb3: num[7:0] = 8'h45;
	8'hb4: num[7:0] = 8'hde;
	8'hb5: num[7:0] = 8'hfd;
	8'hb6: num[7:0] = 8'h8e;
	8'hb7: num[7:0] = 8'h2f;
	8'hb8: num[7:0] = 8'h03;
	8'hb9: num[7:0] = 8'hff;
	8'hba: num[7:0] = 8'h6a;
	8'hbb: num[7:0] = 8'h72;
	8'hbc: num[7:0] = 8'h6d;
	8'hbd: num[7:0] = 8'h6c;
	8'hbe: num[7:0] = 8'h5b;
	8'hbf: num[7:0] = 8'h51;
	8'hc0: num[7:0] = 8'h8d;
	8'hc1: num[7:0] = 8'h1b;
	8'hc2: num[7:0] = 8'haf;
	8'hc3: num[7:0] = 8'h92;
	8'hc4: num[7:0] = 8'hbb;
	8'hc5: num[7:0] = 8'hdd;
	8'hc6: num[7:0] = 8'hbc;
	8'hc7: num[7:0] = 8'h7f;
	8'hc8: num[7:0] = 8'h11;
	8'hc9: num[7:0] = 8'hd9;
	8'hca: num[7:0] = 8'h5c;
	8'hcb: num[7:0] = 8'h41;
	8'hcc: num[7:0] = 8'h1f;
	8'hcd: num[7:0] = 8'h10;
	8'hce: num[7:0] = 8'h5a;
	8'hcf: num[7:0] = 8'hd8;
	8'hd0: num[7:0] = 8'h0a;
	8'hd1: num[7:0] = 8'hc1;
	8'hd2: num[7:0] = 8'h31;
	8'hd3: num[7:0] = 8'h88;
	8'hd4: num[7:0] = 8'ha5;
	8'hd5: num[7:0] = 8'hcd;
	8'hd6: num[7:0] = 8'h7b;
	8'hd7: num[7:0] = 8'hbd;
	8'hd8: num[7:0] = 8'h2d;
	8'hd9: num[7:0] = 8'h74;
	8'hda: num[7:0] = 8'hd0;
	8'hdb: num[7:0] = 8'h12;
	8'hdc: num[7:0] = 8'hb8;
	8'hdd: num[7:0] = 8'he5;
	8'hde: num[7:0] = 8'hb4;
	8'hdf: num[7:0] = 8'hb0;
	8'he0: num[7:0] = 8'h89;
	8'he1: num[7:0] = 8'h69;
	8'he2: num[7:0] = 8'h97;
	8'he3: num[7:0] = 8'h4a;
	8'he4: num[7:0] = 8'h0c;
	8'he5: num[7:0] = 8'h96;
	8'he6: num[7:0] = 8'h77;
	8'he7: num[7:0] = 8'h7e;
	8'he8: num[7:0] = 8'h65;
	8'he9: num[7:0] = 8'hb9;
	8'hea: num[7:0] = 8'hf1;
	8'heb: num[7:0] = 8'h09;
	8'hec: num[7:0] = 8'hc5;
	8'hed: num[7:0] = 8'h6e;
	8'hee: num[7:0] = 8'hc6;
	8'hef: num[7:0] = 8'h84;
	8'hf0: num[7:0] = 8'h18;
	8'hf1: num[7:0] = 8'hf0;
	8'hf2: num[7:0] = 8'h7d;
	8'hf3: num[7:0] = 8'hec;
	8'hf4: num[7:0] = 8'h3a;
	8'hf5: num[7:0] = 8'hdc;
	8'hf6: num[7:0] = 8'h4d;
	8'hf7: num[7:0] = 8'h20;
	8'hf8: num[7:0] = 8'h79;
	8'hf9: num[7:0] = 8'hee;
	8'hfa: num[7:0] = 8'h5f;
	8'hfb: num[7:0] = 8'h3e;
	8'hfc: num[7:0] = 8'hd7;
	8'hfd: num[7:0] = 8'hcb;
	8'hfe: num[7:0] = 8'h39;
	8'hff: num[7:0] = 8'h48;
	default: num[7:0] = 8'h00;
	endcase
	case(num[15:8])
	8'h00: num[15:8] = 8'hd6;
	8'h01: num[15:8] = 8'h90;
	8'h02: num[15:8] = 8'he9;
	8'h03: num[15:8] = 8'hfe;
	8'h04: num[15:8] = 8'hcc;
	8'h05: num[15:8] = 8'he1;
	8'h06: num[15:8] = 8'h3d;
	8'h07: num[15:8] = 8'hb7;
	8'h08: num[15:8] = 8'h16;
	8'h09: num[15:8] = 8'hb6;
	8'h0a: num[15:8] = 8'h14;
	8'h0b: num[15:8] = 8'hc2;
	8'h0c: num[15:8] = 8'h28;
	8'h0d: num[15:8] = 8'hfb;
	8'h0e: num[15:8] = 8'h2c;
	8'h0f: num[15:8] = 8'h05;
	8'h10: num[15:8] = 8'h2b;
	8'h11: num[15:8] = 8'h67;
	8'h12: num[15:8] = 8'h9a;
	8'h13: num[15:8] = 8'h76;
	8'h14: num[15:8] = 8'h2a;
	8'h15: num[15:8] = 8'hbe;
	8'h16: num[15:8] = 8'h04;
	8'h17: num[15:8] = 8'hc3;
	8'h18: num[15:8] = 8'haa;
	8'h19: num[15:8] = 8'h44;
	8'h1a: num[15:8] = 8'h13;
	8'h1b: num[15:8] = 8'h26;
	8'h1c: num[15:8] = 8'h49;
	8'h1d: num[15:8] = 8'h86;
	8'h1e: num[15:8] = 8'h06;
	8'h1f: num[15:8] = 8'h99;
	8'h20: num[15:8] = 8'h9c;
	8'h21: num[15:8] = 8'h42;
	8'h22: num[15:8] = 8'h50;
	8'h23: num[15:8] = 8'hf4;
	8'h24: num[15:8] = 8'h91;
	8'h25: num[15:8] = 8'hef;
	8'h26: num[15:8] = 8'h98;
	8'h27: num[15:8] = 8'h7a;
	8'h28: num[15:8] = 8'h33;
	8'h29: num[15:8] = 8'h54;
	8'h2a: num[15:8] = 8'h0b;
	8'h2b: num[15:8] = 8'h43;
	8'h2c: num[15:8] = 8'hed;
	8'h2d: num[15:8] = 8'hcf;
	8'h2e: num[15:8] = 8'hac;
	8'h2f: num[15:8] = 8'h62;
	8'h30: num[15:8] = 8'he4;
	8'h31: num[15:8] = 8'hb3;
	8'h32: num[15:8] = 8'h1c;
	8'h33: num[15:8] = 8'ha9;
	8'h34: num[15:8] = 8'hc9;
	8'h35: num[15:8] = 8'h08;
	8'h36: num[15:8] = 8'he8;
	8'h37: num[15:8] = 8'h95;
	8'h38: num[15:8] = 8'h80;
	8'h39: num[15:8] = 8'hdf;
	8'h3a: num[15:8] = 8'h94;
	8'h3b: num[15:8] = 8'hfa;
	8'h3c: num[15:8] = 8'h75;
	8'h3d: num[15:8] = 8'h8f;
	8'h3e: num[15:8] = 8'h3f;
	8'h3f: num[15:8] = 8'ha6;
	8'h40: num[15:8] = 8'h47;
	8'h41: num[15:8] = 8'h07;
	8'h42: num[15:8] = 8'ha7;
	8'h43: num[15:8] = 8'hfc;
	8'h44: num[15:8] = 8'hf3;
	8'h45: num[15:8] = 8'h73;
	8'h46: num[15:8] = 8'h17;
	8'h47: num[15:8] = 8'hba;
	8'h48: num[15:8] = 8'h83;
	8'h49: num[15:8] = 8'h59;
	8'h4a: num[15:8] = 8'h3c;
	8'h4b: num[15:8] = 8'h19;
	8'h4c: num[15:8] = 8'he6;
	8'h4d: num[15:8] = 8'h85;
	8'h4e: num[15:8] = 8'h4f;
	8'h4f: num[15:8] = 8'ha8;
	8'h50: num[15:8] = 8'h68;
	8'h51: num[15:8] = 8'h6b;
	8'h52: num[15:8] = 8'h81;
	8'h53: num[15:8] = 8'hb2;
	8'h54: num[15:8] = 8'h71;
	8'h55: num[15:8] = 8'h64;
	8'h56: num[15:8] = 8'hda;
	8'h57: num[15:8] = 8'h8b;
	8'h58: num[15:8] = 8'hf8;
	8'h59: num[15:8] = 8'heb;
	8'h5a: num[15:8] = 8'h0f;
	8'h5b: num[15:8] = 8'h4b;
	8'h5c: num[15:8] = 8'h70;
	8'h5d: num[15:8] = 8'h56;
	8'h5e: num[15:8] = 8'h9d;
	8'h5f: num[15:8] = 8'h35;
	8'h60: num[15:8] = 8'h1e;
	8'h61: num[15:8] = 8'h24;
	8'h62: num[15:8] = 8'h0e;
	8'h63: num[15:8] = 8'h5e;
	8'h64: num[15:8] = 8'h63;
	8'h65: num[15:8] = 8'h58;
	8'h66: num[15:8] = 8'hd1;
	8'h67: num[15:8] = 8'ha2;
	8'h68: num[15:8] = 8'h25;
	8'h69: num[15:8] = 8'h22;
	8'h6a: num[15:8] = 8'h7c;
	8'h6b: num[15:8] = 8'h3b;
	8'h6c: num[15:8] = 8'h01;
	8'h6d: num[15:8] = 8'h21;
	8'h6e: num[15:8] = 8'h78;
	8'h6f: num[15:8] = 8'h87;
	8'h70: num[15:8] = 8'hd4;
	8'h71: num[15:8] = 8'h00;
	8'h72: num[15:8] = 8'h46;
	8'h73: num[15:8] = 8'h57;
	8'h74: num[15:8] = 8'h9f;
	8'h75: num[15:8] = 8'hd3;
	8'h76: num[15:8] = 8'h27;
	8'h77: num[15:8] = 8'h52;
	8'h78: num[15:8] = 8'h4c;
	8'h79: num[15:8] = 8'h36;
	8'h7a: num[15:8] = 8'h02;
	8'h7b: num[15:8] = 8'he7;
	8'h7c: num[15:8] = 8'ha0;
	8'h7d: num[15:8] = 8'hc4;
	8'h7e: num[15:8] = 8'hc8;
	8'h7f: num[15:8] = 8'h9e;
	8'h80: num[15:8] = 8'hea;
	8'h81: num[15:8] = 8'hbf;
	8'h82: num[15:8] = 8'h8a;
	8'h83: num[15:8] = 8'hd2;
	8'h84: num[15:8] = 8'h40;
	8'h85: num[15:8] = 8'hc7;
	8'h86: num[15:8] = 8'h38;
	8'h87: num[15:8] = 8'hb5;
	8'h88: num[15:8] = 8'ha3;
	8'h89: num[15:8] = 8'hf7;
	8'h8a: num[15:8] = 8'hf2;
	8'h8b: num[15:8] = 8'hce;
	8'h8c: num[15:8] = 8'hf9;
	8'h8d: num[15:8] = 8'h61;
	8'h8e: num[15:8] = 8'h15;
	8'h8f: num[15:8] = 8'ha1;
	8'h90: num[15:8] = 8'he0;
	8'h91: num[15:8] = 8'hae;
	8'h92: num[15:8] = 8'h5d;
	8'h93: num[15:8] = 8'ha4;
	8'h94: num[15:8] = 8'h9b;
	8'h95: num[15:8] = 8'h34;
	8'h96: num[15:8] = 8'h1a;
	8'h97: num[15:8] = 8'h55;
	8'h98: num[15:8] = 8'had;
	8'h99: num[15:8] = 8'h93;
	8'h9a: num[15:8] = 8'h32;
	8'h9b: num[15:8] = 8'h30;
	8'h9c: num[15:8] = 8'hf5;
	8'h9d: num[15:8] = 8'h8c;
	8'h9e: num[15:8] = 8'hb1;
	8'h9f: num[15:8] = 8'he3;
	8'ha0: num[15:8] = 8'h1d;
	8'ha1: num[15:8] = 8'hf6;
	8'ha2: num[15:8] = 8'he2;
	8'ha3: num[15:8] = 8'h2e;
	8'ha4: num[15:8] = 8'h82;
	8'ha5: num[15:8] = 8'h66;
	8'ha6: num[15:8] = 8'hca;
	8'ha7: num[15:8] = 8'h60;
	8'ha8: num[15:8] = 8'hc0;
	8'ha9: num[15:8] = 8'h29;
	8'haa: num[15:8] = 8'h23;
	8'hab: num[15:8] = 8'hab;
	8'hac: num[15:8] = 8'h0d;
	8'had: num[15:8] = 8'h53;
	8'hae: num[15:8] = 8'h4e;
	8'haf: num[15:8] = 8'h6f;
	8'hb0: num[15:8] = 8'hd5;
	8'hb1: num[15:8] = 8'hdb;
	8'hb2: num[15:8] = 8'h37;
	8'hb3: num[15:8] = 8'h45;
	8'hb4: num[15:8] = 8'hde;
	8'hb5: num[15:8] = 8'hfd;
	8'hb6: num[15:8] = 8'h8e;
	8'hb7: num[15:8] = 8'h2f;
	8'hb8: num[15:8] = 8'h03;
	8'hb9: num[15:8] = 8'hff;
	8'hba: num[15:8] = 8'h6a;
	8'hbb: num[15:8] = 8'h72;
	8'hbc: num[15:8] = 8'h6d;
	8'hbd: num[15:8] = 8'h6c;
	8'hbe: num[15:8] = 8'h5b;
	8'hbf: num[15:8] = 8'h51;
	8'hc0: num[15:8] = 8'h8d;
	8'hc1: num[15:8] = 8'h1b;
	8'hc2: num[15:8] = 8'haf;
	8'hc3: num[15:8] = 8'h92;
	8'hc4: num[15:8] = 8'hbb;
	8'hc5: num[15:8] = 8'hdd;
	8'hc6: num[15:8] = 8'hbc;
	8'hc7: num[15:8] = 8'h7f;
	8'hc8: num[15:8] = 8'h11;
	8'hc9: num[15:8] = 8'hd9;
	8'hca: num[15:8] = 8'h5c;
	8'hcb: num[15:8] = 8'h41;
	8'hcc: num[15:8] = 8'h1f;
	8'hcd: num[15:8] = 8'h10;
	8'hce: num[15:8] = 8'h5a;
	8'hcf: num[15:8] = 8'hd8;
	8'hd0: num[15:8] = 8'h0a;
	8'hd1: num[15:8] = 8'hc1;
	8'hd2: num[15:8] = 8'h31;
	8'hd3: num[15:8] = 8'h88;
	8'hd4: num[15:8] = 8'ha5;
	8'hd5: num[15:8] = 8'hcd;
	8'hd6: num[15:8] = 8'h7b;
	8'hd7: num[15:8] = 8'hbd;
	8'hd8: num[15:8] = 8'h2d;
	8'hd9: num[15:8] = 8'h74;
	8'hda: num[15:8] = 8'hd0;
	8'hdb: num[15:8] = 8'h12;
	8'hdc: num[15:8] = 8'hb8;
	8'hdd: num[15:8] = 8'he5;
	8'hde: num[15:8] = 8'hb4;
	8'hdf: num[15:8] = 8'hb0;
	8'he0: num[15:8] = 8'h89;
	8'he1: num[15:8] = 8'h69;
	8'he2: num[15:8] = 8'h97;
	8'he3: num[15:8] = 8'h4a;
	8'he4: num[15:8] = 8'h0c;
	8'he5: num[15:8] = 8'h96;
	8'he6: num[15:8] = 8'h77;
	8'he7: num[15:8] = 8'h7e;
	8'he8: num[15:8] = 8'h65;
	8'he9: num[15:8] = 8'hb9;
	8'hea: num[15:8] = 8'hf1;
	8'heb: num[15:8] = 8'h09;
	8'hec: num[15:8] = 8'hc5;
	8'hed: num[15:8] = 8'h6e;
	8'hee: num[15:8] = 8'hc6;
	8'hef: num[15:8] = 8'h84;
	8'hf0: num[15:8] = 8'h18;
	8'hf1: num[15:8] = 8'hf0;
	8'hf2: num[15:8] = 8'h7d;
	8'hf3: num[15:8] = 8'hec;
	8'hf4: num[15:8] = 8'h3a;
	8'hf5: num[15:8] = 8'hdc;
	8'hf6: num[15:8] = 8'h4d;
	8'hf7: num[15:8] = 8'h20;
	8'hf8: num[15:8] = 8'h79;
	8'hf9: num[15:8] = 8'hee;
	8'hfa: num[15:8] = 8'h5f;
	8'hfb: num[15:8] = 8'h3e;
	8'hfc: num[15:8] = 8'hd7;
	8'hfd: num[15:8] = 8'hcb;
	8'hfe: num[15:8] = 8'h39;
	8'hff: num[15:8] = 8'h48;
	default: num[15:8] = 8'h00;
	endcase
	case(num[23:16])
	8'h00: num[23:16] = 8'hd6;
	8'h01: num[23:16] = 8'h90;
	8'h02: num[23:16] = 8'he9;
	8'h03: num[23:16] = 8'hfe;
	8'h04: num[23:16] = 8'hcc;
	8'h05: num[23:16] = 8'he1;
	8'h06: num[23:16] = 8'h3d;
	8'h07: num[23:16] = 8'hb7;
	8'h08: num[23:16] = 8'h16;
	8'h09: num[23:16] = 8'hb6;
	8'h0a: num[23:16] = 8'h14;
	8'h0b: num[23:16] = 8'hc2;
	8'h0c: num[23:16] = 8'h28;
	8'h0d: num[23:16] = 8'hfb;
	8'h0e: num[23:16] = 8'h2c;
	8'h0f: num[23:16] = 8'h05;
	8'h10: num[23:16] = 8'h2b;
	8'h11: num[23:16] = 8'h67;
	8'h12: num[23:16] = 8'h9a;
	8'h13: num[23:16] = 8'h76;
	8'h14: num[23:16] = 8'h2a;
	8'h15: num[23:16] = 8'hbe;
	8'h16: num[23:16] = 8'h04;
	8'h17: num[23:16] = 8'hc3;
	8'h18: num[23:16] = 8'haa;
	8'h19: num[23:16] = 8'h44;
	8'h1a: num[23:16] = 8'h13;
	8'h1b: num[23:16] = 8'h26;
	8'h1c: num[23:16] = 8'h49;
	8'h1d: num[23:16] = 8'h86;
	8'h1e: num[23:16] = 8'h06;
	8'h1f: num[23:16] = 8'h99;
	8'h20: num[23:16] = 8'h9c;
	8'h21: num[23:16] = 8'h42;
	8'h22: num[23:16] = 8'h50;
	8'h23: num[23:16] = 8'hf4;
	8'h24: num[23:16] = 8'h91;
	8'h25: num[23:16] = 8'hef;
	8'h26: num[23:16] = 8'h98;
	8'h27: num[23:16] = 8'h7a;
	8'h28: num[23:16] = 8'h33;
	8'h29: num[23:16] = 8'h54;
	8'h2a: num[23:16] = 8'h0b;
	8'h2b: num[23:16] = 8'h43;
	8'h2c: num[23:16] = 8'hed;
	8'h2d: num[23:16] = 8'hcf;
	8'h2e: num[23:16] = 8'hac;
	8'h2f: num[23:16] = 8'h62;
	8'h30: num[23:16] = 8'he4;
	8'h31: num[23:16] = 8'hb3;
	8'h32: num[23:16] = 8'h1c;
	8'h33: num[23:16] = 8'ha9;
	8'h34: num[23:16] = 8'hc9;
	8'h35: num[23:16] = 8'h08;
	8'h36: num[23:16] = 8'he8;
	8'h37: num[23:16] = 8'h95;
	8'h38: num[23:16] = 8'h80;
	8'h39: num[23:16] = 8'hdf;
	8'h3a: num[23:16] = 8'h94;
	8'h3b: num[23:16] = 8'hfa;
	8'h3c: num[23:16] = 8'h75;
	8'h3d: num[23:16] = 8'h8f;
	8'h3e: num[23:16] = 8'h3f;
	8'h3f: num[23:16] = 8'ha6;
	8'h40: num[23:16] = 8'h47;
	8'h41: num[23:16] = 8'h07;
	8'h42: num[23:16] = 8'ha7;
	8'h43: num[23:16] = 8'hfc;
	8'h44: num[23:16] = 8'hf3;
	8'h45: num[23:16] = 8'h73;
	8'h46: num[23:16] = 8'h17;
	8'h47: num[23:16] = 8'hba;
	8'h48: num[23:16] = 8'h83;
	8'h49: num[23:16] = 8'h59;
	8'h4a: num[23:16] = 8'h3c;
	8'h4b: num[23:16] = 8'h19;
	8'h4c: num[23:16] = 8'he6;
	8'h4d: num[23:16] = 8'h85;
	8'h4e: num[23:16] = 8'h4f;
	8'h4f: num[23:16] = 8'ha8;
	8'h50: num[23:16] = 8'h68;
	8'h51: num[23:16] = 8'h6b;
	8'h52: num[23:16] = 8'h81;
	8'h53: num[23:16] = 8'hb2;
	8'h54: num[23:16] = 8'h71;
	8'h55: num[23:16] = 8'h64;
	8'h56: num[23:16] = 8'hda;
	8'h57: num[23:16] = 8'h8b;
	8'h58: num[23:16] = 8'hf8;
	8'h59: num[23:16] = 8'heb;
	8'h5a: num[23:16] = 8'h0f;
	8'h5b: num[23:16] = 8'h4b;
	8'h5c: num[23:16] = 8'h70;
	8'h5d: num[23:16] = 8'h56;
	8'h5e: num[23:16] = 8'h9d;
	8'h5f: num[23:16] = 8'h35;
	8'h60: num[23:16] = 8'h1e;
	8'h61: num[23:16] = 8'h24;
	8'h62: num[23:16] = 8'h0e;
	8'h63: num[23:16] = 8'h5e;
	8'h64: num[23:16] = 8'h63;
	8'h65: num[23:16] = 8'h58;
	8'h66: num[23:16] = 8'hd1;
	8'h67: num[23:16] = 8'ha2;
	8'h68: num[23:16] = 8'h25;
	8'h69: num[23:16] = 8'h22;
	8'h6a: num[23:16] = 8'h7c;
	8'h6b: num[23:16] = 8'h3b;
	8'h6c: num[23:16] = 8'h01;
	8'h6d: num[23:16] = 8'h21;
	8'h6e: num[23:16] = 8'h78;
	8'h6f: num[23:16] = 8'h87;
	8'h70: num[23:16] = 8'hd4;
	8'h71: num[23:16] = 8'h00;
	8'h72: num[23:16] = 8'h46;
	8'h73: num[23:16] = 8'h57;
	8'h74: num[23:16] = 8'h9f;
	8'h75: num[23:16] = 8'hd3;
	8'h76: num[23:16] = 8'h27;
	8'h77: num[23:16] = 8'h52;
	8'h78: num[23:16] = 8'h4c;
	8'h79: num[23:16] = 8'h36;
	8'h7a: num[23:16] = 8'h02;
	8'h7b: num[23:16] = 8'he7;
	8'h7c: num[23:16] = 8'ha0;
	8'h7d: num[23:16] = 8'hc4;
	8'h7e: num[23:16] = 8'hc8;
	8'h7f: num[23:16] = 8'h9e;
	8'h80: num[23:16] = 8'hea;
	8'h81: num[23:16] = 8'hbf;
	8'h82: num[23:16] = 8'h8a;
	8'h83: num[23:16] = 8'hd2;
	8'h84: num[23:16] = 8'h40;
	8'h85: num[23:16] = 8'hc7;
	8'h86: num[23:16] = 8'h38;
	8'h87: num[23:16] = 8'hb5;
	8'h88: num[23:16] = 8'ha3;
	8'h89: num[23:16] = 8'hf7;
	8'h8a: num[23:16] = 8'hf2;
	8'h8b: num[23:16] = 8'hce;
	8'h8c: num[23:16] = 8'hf9;
	8'h8d: num[23:16] = 8'h61;
	8'h8e: num[23:16] = 8'h15;
	8'h8f: num[23:16] = 8'ha1;
	8'h90: num[23:16] = 8'he0;
	8'h91: num[23:16] = 8'hae;
	8'h92: num[23:16] = 8'h5d;
	8'h93: num[23:16] = 8'ha4;
	8'h94: num[23:16] = 8'h9b;
	8'h95: num[23:16] = 8'h34;
	8'h96: num[23:16] = 8'h1a;
	8'h97: num[23:16] = 8'h55;
	8'h98: num[23:16] = 8'had;
	8'h99: num[23:16] = 8'h93;
	8'h9a: num[23:16] = 8'h32;
	8'h9b: num[23:16] = 8'h30;
	8'h9c: num[23:16] = 8'hf5;
	8'h9d: num[23:16] = 8'h8c;
	8'h9e: num[23:16] = 8'hb1;
	8'h9f: num[23:16] = 8'he3;
	8'ha0: num[23:16] = 8'h1d;
	8'ha1: num[23:16] = 8'hf6;
	8'ha2: num[23:16] = 8'he2;
	8'ha3: num[23:16] = 8'h2e;
	8'ha4: num[23:16] = 8'h82;
	8'ha5: num[23:16] = 8'h66;
	8'ha6: num[23:16] = 8'hca;
	8'ha7: num[23:16] = 8'h60;
	8'ha8: num[23:16] = 8'hc0;
	8'ha9: num[23:16] = 8'h29;
	8'haa: num[23:16] = 8'h23;
	8'hab: num[23:16] = 8'hab;
	8'hac: num[23:16] = 8'h0d;
	8'had: num[23:16] = 8'h53;
	8'hae: num[23:16] = 8'h4e;
	8'haf: num[23:16] = 8'h6f;
	8'hb0: num[23:16] = 8'hd5;
	8'hb1: num[23:16] = 8'hdb;
	8'hb2: num[23:16] = 8'h37;
	8'hb3: num[23:16] = 8'h45;
	8'hb4: num[23:16] = 8'hde;
	8'hb5: num[23:16] = 8'hfd;
	8'hb6: num[23:16] = 8'h8e;
	8'hb7: num[23:16] = 8'h2f;
	8'hb8: num[23:16] = 8'h03;
	8'hb9: num[23:16] = 8'hff;
	8'hba: num[23:16] = 8'h6a;
	8'hbb: num[23:16] = 8'h72;
	8'hbc: num[23:16] = 8'h6d;
	8'hbd: num[23:16] = 8'h6c;
	8'hbe: num[23:16] = 8'h5b;
	8'hbf: num[23:16] = 8'h51;
	8'hc0: num[23:16] = 8'h8d;
	8'hc1: num[23:16] = 8'h1b;
	8'hc2: num[23:16] = 8'haf;
	8'hc3: num[23:16] = 8'h92;
	8'hc4: num[23:16] = 8'hbb;
	8'hc5: num[23:16] = 8'hdd;
	8'hc6: num[23:16] = 8'hbc;
	8'hc7: num[23:16] = 8'h7f;
	8'hc8: num[23:16] = 8'h11;
	8'hc9: num[23:16] = 8'hd9;
	8'hca: num[23:16] = 8'h5c;
	8'hcb: num[23:16] = 8'h41;
	8'hcc: num[23:16] = 8'h1f;
	8'hcd: num[23:16] = 8'h10;
	8'hce: num[23:16] = 8'h5a;
	8'hcf: num[23:16] = 8'hd8;
	8'hd0: num[23:16] = 8'h0a;
	8'hd1: num[23:16] = 8'hc1;
	8'hd2: num[23:16] = 8'h31;
	8'hd3: num[23:16] = 8'h88;
	8'hd4: num[23:16] = 8'ha5;
	8'hd5: num[23:16] = 8'hcd;
	8'hd6: num[23:16] = 8'h7b;
	8'hd7: num[23:16] = 8'hbd;
	8'hd8: num[23:16] = 8'h2d;
	8'hd9: num[23:16] = 8'h74;
	8'hda: num[23:16] = 8'hd0;
	8'hdb: num[23:16] = 8'h12;
	8'hdc: num[23:16] = 8'hb8;
	8'hdd: num[23:16] = 8'he5;
	8'hde: num[23:16] = 8'hb4;
	8'hdf: num[23:16] = 8'hb0;
	8'he0: num[23:16] = 8'h89;
	8'he1: num[23:16] = 8'h69;
	8'he2: num[23:16] = 8'h97;
	8'he3: num[23:16] = 8'h4a;
	8'he4: num[23:16] = 8'h0c;
	8'he5: num[23:16] = 8'h96;
	8'he6: num[23:16] = 8'h77;
	8'he7: num[23:16] = 8'h7e;
	8'he8: num[23:16] = 8'h65;
	8'he9: num[23:16] = 8'hb9;
	8'hea: num[23:16] = 8'hf1;
	8'heb: num[23:16] = 8'h09;
	8'hec: num[23:16] = 8'hc5;
	8'hed: num[23:16] = 8'h6e;
	8'hee: num[23:16] = 8'hc6;
	8'hef: num[23:16] = 8'h84;
	8'hf0: num[23:16] = 8'h18;
	8'hf1: num[23:16] = 8'hf0;
	8'hf2: num[23:16] = 8'h7d;
	8'hf3: num[23:16] = 8'hec;
	8'hf4: num[23:16] = 8'h3a;
	8'hf5: num[23:16] = 8'hdc;
	8'hf6: num[23:16] = 8'h4d;
	8'hf7: num[23:16] = 8'h20;
	8'hf8: num[23:16] = 8'h79;
	8'hf9: num[23:16] = 8'hee;
	8'hfa: num[23:16] = 8'h5f;
	8'hfb: num[23:16] = 8'h3e;
	8'hfc: num[23:16] = 8'hd7;
	8'hfd: num[23:16] = 8'hcb;
	8'hfe: num[23:16] = 8'h39;
	8'hff: num[23:16] = 8'h48;
	default: num[23:16] = 8'h00;
	endcase
	case(num[31:24])
	8'h00: num[31:24] = 8'hd6;
	8'h01: num[31:24] = 8'h90;
	8'h02: num[31:24] = 8'he9;
	8'h03: num[31:24] = 8'hfe;
	8'h04: num[31:24] = 8'hcc;
	8'h05: num[31:24] = 8'he1;
	8'h06: num[31:24] = 8'h3d;
	8'h07: num[31:24] = 8'hb7;
	8'h08: num[31:24] = 8'h16;
	8'h09: num[31:24] = 8'hb6;
	8'h0a: num[31:24] = 8'h14;
	8'h0b: num[31:24] = 8'hc2;
	8'h0c: num[31:24] = 8'h28;
	8'h0d: num[31:24] = 8'hfb;
	8'h0e: num[31:24] = 8'h2c;
	8'h0f: num[31:24] = 8'h05;
	8'h10: num[31:24] = 8'h2b;
	8'h11: num[31:24] = 8'h67;
	8'h12: num[31:24] = 8'h9a;
	8'h13: num[31:24] = 8'h76;
	8'h14: num[31:24] = 8'h2a;
	8'h15: num[31:24] = 8'hbe;
	8'h16: num[31:24] = 8'h04;
	8'h17: num[31:24] = 8'hc3;
	8'h18: num[31:24] = 8'haa;
	8'h19: num[31:24] = 8'h44;
	8'h1a: num[31:24] = 8'h13;
	8'h1b: num[31:24] = 8'h26;
	8'h1c: num[31:24] = 8'h49;
	8'h1d: num[31:24] = 8'h86;
	8'h1e: num[31:24] = 8'h06;
	8'h1f: num[31:24] = 8'h99;
	8'h20: num[31:24] = 8'h9c;
	8'h21: num[31:24] = 8'h42;
	8'h22: num[31:24] = 8'h50;
	8'h23: num[31:24] = 8'hf4;
	8'h24: num[31:24] = 8'h91;
	8'h25: num[31:24] = 8'hef;
	8'h26: num[31:24] = 8'h98;
	8'h27: num[31:24] = 8'h7a;
	8'h28: num[31:24] = 8'h33;
	8'h29: num[31:24] = 8'h54;
	8'h2a: num[31:24] = 8'h0b;
	8'h2b: num[31:24] = 8'h43;
	8'h2c: num[31:24] = 8'hed;
	8'h2d: num[31:24] = 8'hcf;
	8'h2e: num[31:24] = 8'hac;
	8'h2f: num[31:24] = 8'h62;
	8'h30: num[31:24] = 8'he4;
	8'h31: num[31:24] = 8'hb3;
	8'h32: num[31:24] = 8'h1c;
	8'h33: num[31:24] = 8'ha9;
	8'h34: num[31:24] = 8'hc9;
	8'h35: num[31:24] = 8'h08;
	8'h36: num[31:24] = 8'he8;
	8'h37: num[31:24] = 8'h95;
	8'h38: num[31:24] = 8'h80;
	8'h39: num[31:24] = 8'hdf;
	8'h3a: num[31:24] = 8'h94;
	8'h3b: num[31:24] = 8'hfa;
	8'h3c: num[31:24] = 8'h75;
	8'h3d: num[31:24] = 8'h8f;
	8'h3e: num[31:24] = 8'h3f;
	8'h3f: num[31:24] = 8'ha6;
	8'h40: num[31:24] = 8'h47;
	8'h41: num[31:24] = 8'h07;
	8'h42: num[31:24] = 8'ha7;
	8'h43: num[31:24] = 8'hfc;
	8'h44: num[31:24] = 8'hf3;
	8'h45: num[31:24] = 8'h73;
	8'h46: num[31:24] = 8'h17;
	8'h47: num[31:24] = 8'hba;
	8'h48: num[31:24] = 8'h83;
	8'h49: num[31:24] = 8'h59;
	8'h4a: num[31:24] = 8'h3c;
	8'h4b: num[31:24] = 8'h19;
	8'h4c: num[31:24] = 8'he6;
	8'h4d: num[31:24] = 8'h85;
	8'h4e: num[31:24] = 8'h4f;
	8'h4f: num[31:24] = 8'ha8;
	8'h50: num[31:24] = 8'h68;
	8'h51: num[31:24] = 8'h6b;
	8'h52: num[31:24] = 8'h81;
	8'h53: num[31:24] = 8'hb2;
	8'h54: num[31:24] = 8'h71;
	8'h55: num[31:24] = 8'h64;
	8'h56: num[31:24] = 8'hda;
	8'h57: num[31:24] = 8'h8b;
	8'h58: num[31:24] = 8'hf8;
	8'h59: num[31:24] = 8'heb;
	8'h5a: num[31:24] = 8'h0f;
	8'h5b: num[31:24] = 8'h4b;
	8'h5c: num[31:24] = 8'h70;
	8'h5d: num[31:24] = 8'h56;
	8'h5e: num[31:24] = 8'h9d;
	8'h5f: num[31:24] = 8'h35;
	8'h60: num[31:24] = 8'h1e;
	8'h61: num[31:24] = 8'h24;
	8'h62: num[31:24] = 8'h0e;
	8'h63: num[31:24] = 8'h5e;
	8'h64: num[31:24] = 8'h63;
	8'h65: num[31:24] = 8'h58;
	8'h66: num[31:24] = 8'hd1;
	8'h67: num[31:24] = 8'ha2;
	8'h68: num[31:24] = 8'h25;
	8'h69: num[31:24] = 8'h22;
	8'h6a: num[31:24] = 8'h7c;
	8'h6b: num[31:24] = 8'h3b;
	8'h6c: num[31:24] = 8'h01;
	8'h6d: num[31:24] = 8'h21;
	8'h6e: num[31:24] = 8'h78;
	8'h6f: num[31:24] = 8'h87;
	8'h70: num[31:24] = 8'hd4;
	8'h71: num[31:24] = 8'h00;
	8'h72: num[31:24] = 8'h46;
	8'h73: num[31:24] = 8'h57;
	8'h74: num[31:24] = 8'h9f;
	8'h75: num[31:24] = 8'hd3;
	8'h76: num[31:24] = 8'h27;
	8'h77: num[31:24] = 8'h52;
	8'h78: num[31:24] = 8'h4c;
	8'h79: num[31:24] = 8'h36;
	8'h7a: num[31:24] = 8'h02;
	8'h7b: num[31:24] = 8'he7;
	8'h7c: num[31:24] = 8'ha0;
	8'h7d: num[31:24] = 8'hc4;
	8'h7e: num[31:24] = 8'hc8;
	8'h7f: num[31:24] = 8'h9e;
	8'h80: num[31:24] = 8'hea;
	8'h81: num[31:24] = 8'hbf;
	8'h82: num[31:24] = 8'h8a;
	8'h83: num[31:24] = 8'hd2;
	8'h84: num[31:24] = 8'h40;
	8'h85: num[31:24] = 8'hc7;
	8'h86: num[31:24] = 8'h38;
	8'h87: num[31:24] = 8'hb5;
	8'h88: num[31:24] = 8'ha3;
	8'h89: num[31:24] = 8'hf7;
	8'h8a: num[31:24] = 8'hf2;
	8'h8b: num[31:24] = 8'hce;
	8'h8c: num[31:24] = 8'hf9;
	8'h8d: num[31:24] = 8'h61;
	8'h8e: num[31:24] = 8'h15;
	8'h8f: num[31:24] = 8'ha1;
	8'h90: num[31:24] = 8'he0;
	8'h91: num[31:24] = 8'hae;
	8'h92: num[31:24] = 8'h5d;
	8'h93: num[31:24] = 8'ha4;
	8'h94: num[31:24] = 8'h9b;
	8'h95: num[31:24] = 8'h34;
	8'h96: num[31:24] = 8'h1a;
	8'h97: num[31:24] = 8'h55;
	8'h98: num[31:24] = 8'had;
	8'h99: num[31:24] = 8'h93;
	8'h9a: num[31:24] = 8'h32;
	8'h9b: num[31:24] = 8'h30;
	8'h9c: num[31:24] = 8'hf5;
	8'h9d: num[31:24] = 8'h8c;
	8'h9e: num[31:24] = 8'hb1;
	8'h9f: num[31:24] = 8'he3;
	8'ha0: num[31:24] = 8'h1d;
	8'ha1: num[31:24] = 8'hf6;
	8'ha2: num[31:24] = 8'he2;
	8'ha3: num[31:24] = 8'h2e;
	8'ha4: num[31:24] = 8'h82;
	8'ha5: num[31:24] = 8'h66;
	8'ha6: num[31:24] = 8'hca;
	8'ha7: num[31:24] = 8'h60;
	8'ha8: num[31:24] = 8'hc0;
	8'ha9: num[31:24] = 8'h29;
	8'haa: num[31:24] = 8'h23;
	8'hab: num[31:24] = 8'hab;
	8'hac: num[31:24] = 8'h0d;
	8'had: num[31:24] = 8'h53;
	8'hae: num[31:24] = 8'h4e;
	8'haf: num[31:24] = 8'h6f;
	8'hb0: num[31:24] = 8'hd5;
	8'hb1: num[31:24] = 8'hdb;
	8'hb2: num[31:24] = 8'h37;
	8'hb3: num[31:24] = 8'h45;
	8'hb4: num[31:24] = 8'hde;
	8'hb5: num[31:24] = 8'hfd;
	8'hb6: num[31:24] = 8'h8e;
	8'hb7: num[31:24] = 8'h2f;
	8'hb8: num[31:24] = 8'h03;
	8'hb9: num[31:24] = 8'hff;
	8'hba: num[31:24] = 8'h6a;
	8'hbb: num[31:24] = 8'h72;
	8'hbc: num[31:24] = 8'h6d;
	8'hbd: num[31:24] = 8'h6c;
	8'hbe: num[31:24] = 8'h5b;
	8'hbf: num[31:24] = 8'h51;
	8'hc0: num[31:24] = 8'h8d;
	8'hc1: num[31:24] = 8'h1b;
	8'hc2: num[31:24] = 8'haf;
	8'hc3: num[31:24] = 8'h92;
	8'hc4: num[31:24] = 8'hbb;
	8'hc5: num[31:24] = 8'hdd;
	8'hc6: num[31:24] = 8'hbc;
	8'hc7: num[31:24] = 8'h7f;
	8'hc8: num[31:24] = 8'h11;
	8'hc9: num[31:24] = 8'hd9;
	8'hca: num[31:24] = 8'h5c;
	8'hcb: num[31:24] = 8'h41;
	8'hcc: num[31:24] = 8'h1f;
	8'hcd: num[31:24] = 8'h10;
	8'hce: num[31:24] = 8'h5a;
	8'hcf: num[31:24] = 8'hd8;
	8'hd0: num[31:24] = 8'h0a;
	8'hd1: num[31:24] = 8'hc1;
	8'hd2: num[31:24] = 8'h31;
	8'hd3: num[31:24] = 8'h88;
	8'hd4: num[31:24] = 8'ha5;
	8'hd5: num[31:24] = 8'hcd;
	8'hd6: num[31:24] = 8'h7b;
	8'hd7: num[31:24] = 8'hbd;
	8'hd8: num[31:24] = 8'h2d;
	8'hd9: num[31:24] = 8'h74;
	8'hda: num[31:24] = 8'hd0;
	8'hdb: num[31:24] = 8'h12;
	8'hdc: num[31:24] = 8'hb8;
	8'hdd: num[31:24] = 8'he5;
	8'hde: num[31:24] = 8'hb4;
	8'hdf: num[31:24] = 8'hb0;
	8'he0: num[31:24] = 8'h89;
	8'he1: num[31:24] = 8'h69;
	8'he2: num[31:24] = 8'h97;
	8'he3: num[31:24] = 8'h4a;
	8'he4: num[31:24] = 8'h0c;
	8'he5: num[31:24] = 8'h96;
	8'he6: num[31:24] = 8'h77;
	8'he7: num[31:24] = 8'h7e;
	8'he8: num[31:24] = 8'h65;
	8'he9: num[31:24] = 8'hb9;
	8'hea: num[31:24] = 8'hf1;
	8'heb: num[31:24] = 8'h09;
	8'hec: num[31:24] = 8'hc5;
	8'hed: num[31:24] = 8'h6e;
	8'hee: num[31:24] = 8'hc6;
	8'hef: num[31:24] = 8'h84;
	8'hf0: num[31:24] = 8'h18;
	8'hf1: num[31:24] = 8'hf0;
	8'hf2: num[31:24] = 8'h7d;
	8'hf3: num[31:24] = 8'hec;
	8'hf4: num[31:24] = 8'h3a;
	8'hf5: num[31:24] = 8'hdc;
	8'hf6: num[31:24] = 8'h4d;
	8'hf7: num[31:24] = 8'h20;
	8'hf8: num[31:24] = 8'h79;
	8'hf9: num[31:24] = 8'hee;
	8'hfa: num[31:24] = 8'h5f;
	8'hfb: num[31:24] = 8'h3e;
	8'hfc: num[31:24] = 8'hd7;
	8'hfd: num[31:24] = 8'hcb;
	8'hfe: num[31:24] = 8'h39;
	8'hff: num[31:24] = 8'h48;
	default: num[31:24] = 8'h00;
	endcase
        
        RK[i+4] = RK[i] ^ num ^ {num[18:0], num[31:19]} ^ {num[8:0], num[31:9]};
    end
   
    
    text[0] = plain[127:96];
    text[1] = plain[95:64];
    text[2] = plain[63:32];
    text[3] = plain[31:0];  
    for(i = 0; i < 32; i = i + 1)begin
        num = text[i+1] ^ text[i+2] ^text[i+3] ^ RK[i+4];
        
    case(num[7:0])
	8'h00: num[7:0] = 8'hd6;
	8'h01: num[7:0] = 8'h90;
	8'h02: num[7:0] = 8'he9;
	8'h03: num[7:0] = 8'hfe;
	8'h04: num[7:0] = 8'hcc;
	8'h05: num[7:0] = 8'he1;
	8'h06: num[7:0] = 8'h3d;
	8'h07: num[7:0] = 8'hb7;
	8'h08: num[7:0] = 8'h16;
	8'h09: num[7:0] = 8'hb6;
	8'h0a: num[7:0] = 8'h14;
	8'h0b: num[7:0] = 8'hc2;
	8'h0c: num[7:0] = 8'h28;
	8'h0d: num[7:0] = 8'hfb;
	8'h0e: num[7:0] = 8'h2c;
	8'h0f: num[7:0] = 8'h05;
	8'h10: num[7:0] = 8'h2b;
	8'h11: num[7:0] = 8'h67;
	8'h12: num[7:0] = 8'h9a;
	8'h13: num[7:0] = 8'h76;
	8'h14: num[7:0] = 8'h2a;
	8'h15: num[7:0] = 8'hbe;
	8'h16: num[7:0] = 8'h04;
	8'h17: num[7:0] = 8'hc3;
	8'h18: num[7:0] = 8'haa;
	8'h19: num[7:0] = 8'h44;
	8'h1a: num[7:0] = 8'h13;
	8'h1b: num[7:0] = 8'h26;
	8'h1c: num[7:0] = 8'h49;
	8'h1d: num[7:0] = 8'h86;
	8'h1e: num[7:0] = 8'h06;
	8'h1f: num[7:0] = 8'h99;
	8'h20: num[7:0] = 8'h9c;
	8'h21: num[7:0] = 8'h42;
	8'h22: num[7:0] = 8'h50;
	8'h23: num[7:0] = 8'hf4;
	8'h24: num[7:0] = 8'h91;
	8'h25: num[7:0] = 8'hef;
	8'h26: num[7:0] = 8'h98;
	8'h27: num[7:0] = 8'h7a;
	8'h28: num[7:0] = 8'h33;
	8'h29: num[7:0] = 8'h54;
	8'h2a: num[7:0] = 8'h0b;
	8'h2b: num[7:0] = 8'h43;
	8'h2c: num[7:0] = 8'hed;
	8'h2d: num[7:0] = 8'hcf;
	8'h2e: num[7:0] = 8'hac;
	8'h2f: num[7:0] = 8'h62;
	8'h30: num[7:0] = 8'he4;
	8'h31: num[7:0] = 8'hb3;
	8'h32: num[7:0] = 8'h1c;
	8'h33: num[7:0] = 8'ha9;
	8'h34: num[7:0] = 8'hc9;
	8'h35: num[7:0] = 8'h08;
	8'h36: num[7:0] = 8'he8;
	8'h37: num[7:0] = 8'h95;
	8'h38: num[7:0] = 8'h80;
	8'h39: num[7:0] = 8'hdf;
	8'h3a: num[7:0] = 8'h94;
	8'h3b: num[7:0] = 8'hfa;
	8'h3c: num[7:0] = 8'h75;
	8'h3d: num[7:0] = 8'h8f;
	8'h3e: num[7:0] = 8'h3f;
	8'h3f: num[7:0] = 8'ha6;
	8'h40: num[7:0] = 8'h47;
	8'h41: num[7:0] = 8'h07;
	8'h42: num[7:0] = 8'ha7;
	8'h43: num[7:0] = 8'hfc;
	8'h44: num[7:0] = 8'hf3;
	8'h45: num[7:0] = 8'h73;
	8'h46: num[7:0] = 8'h17;
	8'h47: num[7:0] = 8'hba;
	8'h48: num[7:0] = 8'h83;
	8'h49: num[7:0] = 8'h59;
	8'h4a: num[7:0] = 8'h3c;
	8'h4b: num[7:0] = 8'h19;
	8'h4c: num[7:0] = 8'he6;
	8'h4d: num[7:0] = 8'h85;
	8'h4e: num[7:0] = 8'h4f;
	8'h4f: num[7:0] = 8'ha8;
	8'h50: num[7:0] = 8'h68;
	8'h51: num[7:0] = 8'h6b;
	8'h52: num[7:0] = 8'h81;
	8'h53: num[7:0] = 8'hb2;
	8'h54: num[7:0] = 8'h71;
	8'h55: num[7:0] = 8'h64;
	8'h56: num[7:0] = 8'hda;
	8'h57: num[7:0] = 8'h8b;
	8'h58: num[7:0] = 8'hf8;
	8'h59: num[7:0] = 8'heb;
	8'h5a: num[7:0] = 8'h0f;
	8'h5b: num[7:0] = 8'h4b;
	8'h5c: num[7:0] = 8'h70;
	8'h5d: num[7:0] = 8'h56;
	8'h5e: num[7:0] = 8'h9d;
	8'h5f: num[7:0] = 8'h35;
	8'h60: num[7:0] = 8'h1e;
	8'h61: num[7:0] = 8'h24;
	8'h62: num[7:0] = 8'h0e;
	8'h63: num[7:0] = 8'h5e;
	8'h64: num[7:0] = 8'h63;
	8'h65: num[7:0] = 8'h58;
	8'h66: num[7:0] = 8'hd1;
	8'h67: num[7:0] = 8'ha2;
	8'h68: num[7:0] = 8'h25;
	8'h69: num[7:0] = 8'h22;
	8'h6a: num[7:0] = 8'h7c;
	8'h6b: num[7:0] = 8'h3b;
	8'h6c: num[7:0] = 8'h01;
	8'h6d: num[7:0] = 8'h21;
	8'h6e: num[7:0] = 8'h78;
	8'h6f: num[7:0] = 8'h87;
	8'h70: num[7:0] = 8'hd4;
	8'h71: num[7:0] = 8'h00;
	8'h72: num[7:0] = 8'h46;
	8'h73: num[7:0] = 8'h57;
	8'h74: num[7:0] = 8'h9f;
	8'h75: num[7:0] = 8'hd3;
	8'h76: num[7:0] = 8'h27;
	8'h77: num[7:0] = 8'h52;
	8'h78: num[7:0] = 8'h4c;
	8'h79: num[7:0] = 8'h36;
	8'h7a: num[7:0] = 8'h02;
	8'h7b: num[7:0] = 8'he7;
	8'h7c: num[7:0] = 8'ha0;
	8'h7d: num[7:0] = 8'hc4;
	8'h7e: num[7:0] = 8'hc8;
	8'h7f: num[7:0] = 8'h9e;
	8'h80: num[7:0] = 8'hea;
	8'h81: num[7:0] = 8'hbf;
	8'h82: num[7:0] = 8'h8a;
	8'h83: num[7:0] = 8'hd2;
	8'h84: num[7:0] = 8'h40;
	8'h85: num[7:0] = 8'hc7;
	8'h86: num[7:0] = 8'h38;
	8'h87: num[7:0] = 8'hb5;
	8'h88: num[7:0] = 8'ha3;
	8'h89: num[7:0] = 8'hf7;
	8'h8a: num[7:0] = 8'hf2;
	8'h8b: num[7:0] = 8'hce;
	8'h8c: num[7:0] = 8'hf9;
	8'h8d: num[7:0] = 8'h61;
	8'h8e: num[7:0] = 8'h15;
	8'h8f: num[7:0] = 8'ha1;
	8'h90: num[7:0] = 8'he0;
	8'h91: num[7:0] = 8'hae;
	8'h92: num[7:0] = 8'h5d;
	8'h93: num[7:0] = 8'ha4;
	8'h94: num[7:0] = 8'h9b;
	8'h95: num[7:0] = 8'h34;
	8'h96: num[7:0] = 8'h1a;
	8'h97: num[7:0] = 8'h55;
	8'h98: num[7:0] = 8'had;
	8'h99: num[7:0] = 8'h93;
	8'h9a: num[7:0] = 8'h32;
	8'h9b: num[7:0] = 8'h30;
	8'h9c: num[7:0] = 8'hf5;
	8'h9d: num[7:0] = 8'h8c;
	8'h9e: num[7:0] = 8'hb1;
	8'h9f: num[7:0] = 8'he3;
	8'ha0: num[7:0] = 8'h1d;
	8'ha1: num[7:0] = 8'hf6;
	8'ha2: num[7:0] = 8'he2;
	8'ha3: num[7:0] = 8'h2e;
	8'ha4: num[7:0] = 8'h82;
	8'ha5: num[7:0] = 8'h66;
	8'ha6: num[7:0] = 8'hca;
	8'ha7: num[7:0] = 8'h60;
	8'ha8: num[7:0] = 8'hc0;
	8'ha9: num[7:0] = 8'h29;
	8'haa: num[7:0] = 8'h23;
	8'hab: num[7:0] = 8'hab;
	8'hac: num[7:0] = 8'h0d;
	8'had: num[7:0] = 8'h53;
	8'hae: num[7:0] = 8'h4e;
	8'haf: num[7:0] = 8'h6f;
	8'hb0: num[7:0] = 8'hd5;
	8'hb1: num[7:0] = 8'hdb;
	8'hb2: num[7:0] = 8'h37;
	8'hb3: num[7:0] = 8'h45;
	8'hb4: num[7:0] = 8'hde;
	8'hb5: num[7:0] = 8'hfd;
	8'hb6: num[7:0] = 8'h8e;
	8'hb7: num[7:0] = 8'h2f;
	8'hb8: num[7:0] = 8'h03;
	8'hb9: num[7:0] = 8'hff;
	8'hba: num[7:0] = 8'h6a;
	8'hbb: num[7:0] = 8'h72;
	8'hbc: num[7:0] = 8'h6d;
	8'hbd: num[7:0] = 8'h6c;
	8'hbe: num[7:0] = 8'h5b;
	8'hbf: num[7:0] = 8'h51;
	8'hc0: num[7:0] = 8'h8d;
	8'hc1: num[7:0] = 8'h1b;
	8'hc2: num[7:0] = 8'haf;
	8'hc3: num[7:0] = 8'h92;
	8'hc4: num[7:0] = 8'hbb;
	8'hc5: num[7:0] = 8'hdd;
	8'hc6: num[7:0] = 8'hbc;
	8'hc7: num[7:0] = 8'h7f;
	8'hc8: num[7:0] = 8'h11;
	8'hc9: num[7:0] = 8'hd9;
	8'hca: num[7:0] = 8'h5c;
	8'hcb: num[7:0] = 8'h41;
	8'hcc: num[7:0] = 8'h1f;
	8'hcd: num[7:0] = 8'h10;
	8'hce: num[7:0] = 8'h5a;
	8'hcf: num[7:0] = 8'hd8;
	8'hd0: num[7:0] = 8'h0a;
	8'hd1: num[7:0] = 8'hc1;
	8'hd2: num[7:0] = 8'h31;
	8'hd3: num[7:0] = 8'h88;
	8'hd4: num[7:0] = 8'ha5;
	8'hd5: num[7:0] = 8'hcd;
	8'hd6: num[7:0] = 8'h7b;
	8'hd7: num[7:0] = 8'hbd;
	8'hd8: num[7:0] = 8'h2d;
	8'hd9: num[7:0] = 8'h74;
	8'hda: num[7:0] = 8'hd0;
	8'hdb: num[7:0] = 8'h12;
	8'hdc: num[7:0] = 8'hb8;
	8'hdd: num[7:0] = 8'he5;
	8'hde: num[7:0] = 8'hb4;
	8'hdf: num[7:0] = 8'hb0;
	8'he0: num[7:0] = 8'h89;
	8'he1: num[7:0] = 8'h69;
	8'he2: num[7:0] = 8'h97;
	8'he3: num[7:0] = 8'h4a;
	8'he4: num[7:0] = 8'h0c;
	8'he5: num[7:0] = 8'h96;
	8'he6: num[7:0] = 8'h77;
	8'he7: num[7:0] = 8'h7e;
	8'he8: num[7:0] = 8'h65;
	8'he9: num[7:0] = 8'hb9;
	8'hea: num[7:0] = 8'hf1;
	8'heb: num[7:0] = 8'h09;
	8'hec: num[7:0] = 8'hc5;
	8'hed: num[7:0] = 8'h6e;
	8'hee: num[7:0] = 8'hc6;
	8'hef: num[7:0] = 8'h84;
	8'hf0: num[7:0] = 8'h18;
	8'hf1: num[7:0] = 8'hf0;
	8'hf2: num[7:0] = 8'h7d;
	8'hf3: num[7:0] = 8'hec;
	8'hf4: num[7:0] = 8'h3a;
	8'hf5: num[7:0] = 8'hdc;
	8'hf6: num[7:0] = 8'h4d;
	8'hf7: num[7:0] = 8'h20;
	8'hf8: num[7:0] = 8'h79;
	8'hf9: num[7:0] = 8'hee;
	8'hfa: num[7:0] = 8'h5f;
	8'hfb: num[7:0] = 8'h3e;
	8'hfc: num[7:0] = 8'hd7;
	8'hfd: num[7:0] = 8'hcb;
	8'hfe: num[7:0] = 8'h39;
	8'hff: num[7:0] = 8'h48;
	default: num[7:0] = 8'h00;
	endcase
	case(num[15:8])
	8'h00: num[15:8] = 8'hd6;
	8'h01: num[15:8] = 8'h90;
	8'h02: num[15:8] = 8'he9;
	8'h03: num[15:8] = 8'hfe;
	8'h04: num[15:8] = 8'hcc;
	8'h05: num[15:8] = 8'he1;
	8'h06: num[15:8] = 8'h3d;
	8'h07: num[15:8] = 8'hb7;
	8'h08: num[15:8] = 8'h16;
	8'h09: num[15:8] = 8'hb6;
	8'h0a: num[15:8] = 8'h14;
	8'h0b: num[15:8] = 8'hc2;
	8'h0c: num[15:8] = 8'h28;
	8'h0d: num[15:8] = 8'hfb;
	8'h0e: num[15:8] = 8'h2c;
	8'h0f: num[15:8] = 8'h05;
	8'h10: num[15:8] = 8'h2b;
	8'h11: num[15:8] = 8'h67;
	8'h12: num[15:8] = 8'h9a;
	8'h13: num[15:8] = 8'h76;
	8'h14: num[15:8] = 8'h2a;
	8'h15: num[15:8] = 8'hbe;
	8'h16: num[15:8] = 8'h04;
	8'h17: num[15:8] = 8'hc3;
	8'h18: num[15:8] = 8'haa;
	8'h19: num[15:8] = 8'h44;
	8'h1a: num[15:8] = 8'h13;
	8'h1b: num[15:8] = 8'h26;
	8'h1c: num[15:8] = 8'h49;
	8'h1d: num[15:8] = 8'h86;
	8'h1e: num[15:8] = 8'h06;
	8'h1f: num[15:8] = 8'h99;
	8'h20: num[15:8] = 8'h9c;
	8'h21: num[15:8] = 8'h42;
	8'h22: num[15:8] = 8'h50;
	8'h23: num[15:8] = 8'hf4;
	8'h24: num[15:8] = 8'h91;
	8'h25: num[15:8] = 8'hef;
	8'h26: num[15:8] = 8'h98;
	8'h27: num[15:8] = 8'h7a;
	8'h28: num[15:8] = 8'h33;
	8'h29: num[15:8] = 8'h54;
	8'h2a: num[15:8] = 8'h0b;
	8'h2b: num[15:8] = 8'h43;
	8'h2c: num[15:8] = 8'hed;
	8'h2d: num[15:8] = 8'hcf;
	8'h2e: num[15:8] = 8'hac;
	8'h2f: num[15:8] = 8'h62;
	8'h30: num[15:8] = 8'he4;
	8'h31: num[15:8] = 8'hb3;
	8'h32: num[15:8] = 8'h1c;
	8'h33: num[15:8] = 8'ha9;
	8'h34: num[15:8] = 8'hc9;
	8'h35: num[15:8] = 8'h08;
	8'h36: num[15:8] = 8'he8;
	8'h37: num[15:8] = 8'h95;
	8'h38: num[15:8] = 8'h80;
	8'h39: num[15:8] = 8'hdf;
	8'h3a: num[15:8] = 8'h94;
	8'h3b: num[15:8] = 8'hfa;
	8'h3c: num[15:8] = 8'h75;
	8'h3d: num[15:8] = 8'h8f;
	8'h3e: num[15:8] = 8'h3f;
	8'h3f: num[15:8] = 8'ha6;
	8'h40: num[15:8] = 8'h47;
	8'h41: num[15:8] = 8'h07;
	8'h42: num[15:8] = 8'ha7;
	8'h43: num[15:8] = 8'hfc;
	8'h44: num[15:8] = 8'hf3;
	8'h45: num[15:8] = 8'h73;
	8'h46: num[15:8] = 8'h17;
	8'h47: num[15:8] = 8'hba;
	8'h48: num[15:8] = 8'h83;
	8'h49: num[15:8] = 8'h59;
	8'h4a: num[15:8] = 8'h3c;
	8'h4b: num[15:8] = 8'h19;
	8'h4c: num[15:8] = 8'he6;
	8'h4d: num[15:8] = 8'h85;
	8'h4e: num[15:8] = 8'h4f;
	8'h4f: num[15:8] = 8'ha8;
	8'h50: num[15:8] = 8'h68;
	8'h51: num[15:8] = 8'h6b;
	8'h52: num[15:8] = 8'h81;
	8'h53: num[15:8] = 8'hb2;
	8'h54: num[15:8] = 8'h71;
	8'h55: num[15:8] = 8'h64;
	8'h56: num[15:8] = 8'hda;
	8'h57: num[15:8] = 8'h8b;
	8'h58: num[15:8] = 8'hf8;
	8'h59: num[15:8] = 8'heb;
	8'h5a: num[15:8] = 8'h0f;
	8'h5b: num[15:8] = 8'h4b;
	8'h5c: num[15:8] = 8'h70;
	8'h5d: num[15:8] = 8'h56;
	8'h5e: num[15:8] = 8'h9d;
	8'h5f: num[15:8] = 8'h35;
	8'h60: num[15:8] = 8'h1e;
	8'h61: num[15:8] = 8'h24;
	8'h62: num[15:8] = 8'h0e;
	8'h63: num[15:8] = 8'h5e;
	8'h64: num[15:8] = 8'h63;
	8'h65: num[15:8] = 8'h58;
	8'h66: num[15:8] = 8'hd1;
	8'h67: num[15:8] = 8'ha2;
	8'h68: num[15:8] = 8'h25;
	8'h69: num[15:8] = 8'h22;
	8'h6a: num[15:8] = 8'h7c;
	8'h6b: num[15:8] = 8'h3b;
	8'h6c: num[15:8] = 8'h01;
	8'h6d: num[15:8] = 8'h21;
	8'h6e: num[15:8] = 8'h78;
	8'h6f: num[15:8] = 8'h87;
	8'h70: num[15:8] = 8'hd4;
	8'h71: num[15:8] = 8'h00;
	8'h72: num[15:8] = 8'h46;
	8'h73: num[15:8] = 8'h57;
	8'h74: num[15:8] = 8'h9f;
	8'h75: num[15:8] = 8'hd3;
	8'h76: num[15:8] = 8'h27;
	8'h77: num[15:8] = 8'h52;
	8'h78: num[15:8] = 8'h4c;
	8'h79: num[15:8] = 8'h36;
	8'h7a: num[15:8] = 8'h02;
	8'h7b: num[15:8] = 8'he7;
	8'h7c: num[15:8] = 8'ha0;
	8'h7d: num[15:8] = 8'hc4;
	8'h7e: num[15:8] = 8'hc8;
	8'h7f: num[15:8] = 8'h9e;
	8'h80: num[15:8] = 8'hea;
	8'h81: num[15:8] = 8'hbf;
	8'h82: num[15:8] = 8'h8a;
	8'h83: num[15:8] = 8'hd2;
	8'h84: num[15:8] = 8'h40;
	8'h85: num[15:8] = 8'hc7;
	8'h86: num[15:8] = 8'h38;
	8'h87: num[15:8] = 8'hb5;
	8'h88: num[15:8] = 8'ha3;
	8'h89: num[15:8] = 8'hf7;
	8'h8a: num[15:8] = 8'hf2;
	8'h8b: num[15:8] = 8'hce;
	8'h8c: num[15:8] = 8'hf9;
	8'h8d: num[15:8] = 8'h61;
	8'h8e: num[15:8] = 8'h15;
	8'h8f: num[15:8] = 8'ha1;
	8'h90: num[15:8] = 8'he0;
	8'h91: num[15:8] = 8'hae;
	8'h92: num[15:8] = 8'h5d;
	8'h93: num[15:8] = 8'ha4;
	8'h94: num[15:8] = 8'h9b;
	8'h95: num[15:8] = 8'h34;
	8'h96: num[15:8] = 8'h1a;
	8'h97: num[15:8] = 8'h55;
	8'h98: num[15:8] = 8'had;
	8'h99: num[15:8] = 8'h93;
	8'h9a: num[15:8] = 8'h32;
	8'h9b: num[15:8] = 8'h30;
	8'h9c: num[15:8] = 8'hf5;
	8'h9d: num[15:8] = 8'h8c;
	8'h9e: num[15:8] = 8'hb1;
	8'h9f: num[15:8] = 8'he3;
	8'ha0: num[15:8] = 8'h1d;
	8'ha1: num[15:8] = 8'hf6;
	8'ha2: num[15:8] = 8'he2;
	8'ha3: num[15:8] = 8'h2e;
	8'ha4: num[15:8] = 8'h82;
	8'ha5: num[15:8] = 8'h66;
	8'ha6: num[15:8] = 8'hca;
	8'ha7: num[15:8] = 8'h60;
	8'ha8: num[15:8] = 8'hc0;
	8'ha9: num[15:8] = 8'h29;
	8'haa: num[15:8] = 8'h23;
	8'hab: num[15:8] = 8'hab;
	8'hac: num[15:8] = 8'h0d;
	8'had: num[15:8] = 8'h53;
	8'hae: num[15:8] = 8'h4e;
	8'haf: num[15:8] = 8'h6f;
	8'hb0: num[15:8] = 8'hd5;
	8'hb1: num[15:8] = 8'hdb;
	8'hb2: num[15:8] = 8'h37;
	8'hb3: num[15:8] = 8'h45;
	8'hb4: num[15:8] = 8'hde;
	8'hb5: num[15:8] = 8'hfd;
	8'hb6: num[15:8] = 8'h8e;
	8'hb7: num[15:8] = 8'h2f;
	8'hb8: num[15:8] = 8'h03;
	8'hb9: num[15:8] = 8'hff;
	8'hba: num[15:8] = 8'h6a;
	8'hbb: num[15:8] = 8'h72;
	8'hbc: num[15:8] = 8'h6d;
	8'hbd: num[15:8] = 8'h6c;
	8'hbe: num[15:8] = 8'h5b;
	8'hbf: num[15:8] = 8'h51;
	8'hc0: num[15:8] = 8'h8d;
	8'hc1: num[15:8] = 8'h1b;
	8'hc2: num[15:8] = 8'haf;
	8'hc3: num[15:8] = 8'h92;
	8'hc4: num[15:8] = 8'hbb;
	8'hc5: num[15:8] = 8'hdd;
	8'hc6: num[15:8] = 8'hbc;
	8'hc7: num[15:8] = 8'h7f;
	8'hc8: num[15:8] = 8'h11;
	8'hc9: num[15:8] = 8'hd9;
	8'hca: num[15:8] = 8'h5c;
	8'hcb: num[15:8] = 8'h41;
	8'hcc: num[15:8] = 8'h1f;
	8'hcd: num[15:8] = 8'h10;
	8'hce: num[15:8] = 8'h5a;
	8'hcf: num[15:8] = 8'hd8;
	8'hd0: num[15:8] = 8'h0a;
	8'hd1: num[15:8] = 8'hc1;
	8'hd2: num[15:8] = 8'h31;
	8'hd3: num[15:8] = 8'h88;
	8'hd4: num[15:8] = 8'ha5;
	8'hd5: num[15:8] = 8'hcd;
	8'hd6: num[15:8] = 8'h7b;
	8'hd7: num[15:8] = 8'hbd;
	8'hd8: num[15:8] = 8'h2d;
	8'hd9: num[15:8] = 8'h74;
	8'hda: num[15:8] = 8'hd0;
	8'hdb: num[15:8] = 8'h12;
	8'hdc: num[15:8] = 8'hb8;
	8'hdd: num[15:8] = 8'he5;
	8'hde: num[15:8] = 8'hb4;
	8'hdf: num[15:8] = 8'hb0;
	8'he0: num[15:8] = 8'h89;
	8'he1: num[15:8] = 8'h69;
	8'he2: num[15:8] = 8'h97;
	8'he3: num[15:8] = 8'h4a;
	8'he4: num[15:8] = 8'h0c;
	8'he5: num[15:8] = 8'h96;
	8'he6: num[15:8] = 8'h77;
	8'he7: num[15:8] = 8'h7e;
	8'he8: num[15:8] = 8'h65;
	8'he9: num[15:8] = 8'hb9;
	8'hea: num[15:8] = 8'hf1;
	8'heb: num[15:8] = 8'h09;
	8'hec: num[15:8] = 8'hc5;
	8'hed: num[15:8] = 8'h6e;
	8'hee: num[15:8] = 8'hc6;
	8'hef: num[15:8] = 8'h84;
	8'hf0: num[15:8] = 8'h18;
	8'hf1: num[15:8] = 8'hf0;
	8'hf2: num[15:8] = 8'h7d;
	8'hf3: num[15:8] = 8'hec;
	8'hf4: num[15:8] = 8'h3a;
	8'hf5: num[15:8] = 8'hdc;
	8'hf6: num[15:8] = 8'h4d;
	8'hf7: num[15:8] = 8'h20;
	8'hf8: num[15:8] = 8'h79;
	8'hf9: num[15:8] = 8'hee;
	8'hfa: num[15:8] = 8'h5f;
	8'hfb: num[15:8] = 8'h3e;
	8'hfc: num[15:8] = 8'hd7;
	8'hfd: num[15:8] = 8'hcb;
	8'hfe: num[15:8] = 8'h39;
	8'hff: num[15:8] = 8'h48;
	default: num[15:8] = 8'h00;
	endcase
	case(num[23:16])
	8'h00: num[23:16] = 8'hd6;
	8'h01: num[23:16] = 8'h90;
	8'h02: num[23:16] = 8'he9;
	8'h03: num[23:16] = 8'hfe;
	8'h04: num[23:16] = 8'hcc;
	8'h05: num[23:16] = 8'he1;
	8'h06: num[23:16] = 8'h3d;
	8'h07: num[23:16] = 8'hb7;
	8'h08: num[23:16] = 8'h16;
	8'h09: num[23:16] = 8'hb6;
	8'h0a: num[23:16] = 8'h14;
	8'h0b: num[23:16] = 8'hc2;
	8'h0c: num[23:16] = 8'h28;
	8'h0d: num[23:16] = 8'hfb;
	8'h0e: num[23:16] = 8'h2c;
	8'h0f: num[23:16] = 8'h05;
	8'h10: num[23:16] = 8'h2b;
	8'h11: num[23:16] = 8'h67;
	8'h12: num[23:16] = 8'h9a;
	8'h13: num[23:16] = 8'h76;
	8'h14: num[23:16] = 8'h2a;
	8'h15: num[23:16] = 8'hbe;
	8'h16: num[23:16] = 8'h04;
	8'h17: num[23:16] = 8'hc3;
	8'h18: num[23:16] = 8'haa;
	8'h19: num[23:16] = 8'h44;
	8'h1a: num[23:16] = 8'h13;
	8'h1b: num[23:16] = 8'h26;
	8'h1c: num[23:16] = 8'h49;
	8'h1d: num[23:16] = 8'h86;
	8'h1e: num[23:16] = 8'h06;
	8'h1f: num[23:16] = 8'h99;
	8'h20: num[23:16] = 8'h9c;
	8'h21: num[23:16] = 8'h42;
	8'h22: num[23:16] = 8'h50;
	8'h23: num[23:16] = 8'hf4;
	8'h24: num[23:16] = 8'h91;
	8'h25: num[23:16] = 8'hef;
	8'h26: num[23:16] = 8'h98;
	8'h27: num[23:16] = 8'h7a;
	8'h28: num[23:16] = 8'h33;
	8'h29: num[23:16] = 8'h54;
	8'h2a: num[23:16] = 8'h0b;
	8'h2b: num[23:16] = 8'h43;
	8'h2c: num[23:16] = 8'hed;
	8'h2d: num[23:16] = 8'hcf;
	8'h2e: num[23:16] = 8'hac;
	8'h2f: num[23:16] = 8'h62;
	8'h30: num[23:16] = 8'he4;
	8'h31: num[23:16] = 8'hb3;
	8'h32: num[23:16] = 8'h1c;
	8'h33: num[23:16] = 8'ha9;
	8'h34: num[23:16] = 8'hc9;
	8'h35: num[23:16] = 8'h08;
	8'h36: num[23:16] = 8'he8;
	8'h37: num[23:16] = 8'h95;
	8'h38: num[23:16] = 8'h80;
	8'h39: num[23:16] = 8'hdf;
	8'h3a: num[23:16] = 8'h94;
	8'h3b: num[23:16] = 8'hfa;
	8'h3c: num[23:16] = 8'h75;
	8'h3d: num[23:16] = 8'h8f;
	8'h3e: num[23:16] = 8'h3f;
	8'h3f: num[23:16] = 8'ha6;
	8'h40: num[23:16] = 8'h47;
	8'h41: num[23:16] = 8'h07;
	8'h42: num[23:16] = 8'ha7;
	8'h43: num[23:16] = 8'hfc;
	8'h44: num[23:16] = 8'hf3;
	8'h45: num[23:16] = 8'h73;
	8'h46: num[23:16] = 8'h17;
	8'h47: num[23:16] = 8'hba;
	8'h48: num[23:16] = 8'h83;
	8'h49: num[23:16] = 8'h59;
	8'h4a: num[23:16] = 8'h3c;
	8'h4b: num[23:16] = 8'h19;
	8'h4c: num[23:16] = 8'he6;
	8'h4d: num[23:16] = 8'h85;
	8'h4e: num[23:16] = 8'h4f;
	8'h4f: num[23:16] = 8'ha8;
	8'h50: num[23:16] = 8'h68;
	8'h51: num[23:16] = 8'h6b;
	8'h52: num[23:16] = 8'h81;
	8'h53: num[23:16] = 8'hb2;
	8'h54: num[23:16] = 8'h71;
	8'h55: num[23:16] = 8'h64;
	8'h56: num[23:16] = 8'hda;
	8'h57: num[23:16] = 8'h8b;
	8'h58: num[23:16] = 8'hf8;
	8'h59: num[23:16] = 8'heb;
	8'h5a: num[23:16] = 8'h0f;
	8'h5b: num[23:16] = 8'h4b;
	8'h5c: num[23:16] = 8'h70;
	8'h5d: num[23:16] = 8'h56;
	8'h5e: num[23:16] = 8'h9d;
	8'h5f: num[23:16] = 8'h35;
	8'h60: num[23:16] = 8'h1e;
	8'h61: num[23:16] = 8'h24;
	8'h62: num[23:16] = 8'h0e;
	8'h63: num[23:16] = 8'h5e;
	8'h64: num[23:16] = 8'h63;
	8'h65: num[23:16] = 8'h58;
	8'h66: num[23:16] = 8'hd1;
	8'h67: num[23:16] = 8'ha2;
	8'h68: num[23:16] = 8'h25;
	8'h69: num[23:16] = 8'h22;
	8'h6a: num[23:16] = 8'h7c;
	8'h6b: num[23:16] = 8'h3b;
	8'h6c: num[23:16] = 8'h01;
	8'h6d: num[23:16] = 8'h21;
	8'h6e: num[23:16] = 8'h78;
	8'h6f: num[23:16] = 8'h87;
	8'h70: num[23:16] = 8'hd4;
	8'h71: num[23:16] = 8'h00;
	8'h72: num[23:16] = 8'h46;
	8'h73: num[23:16] = 8'h57;
	8'h74: num[23:16] = 8'h9f;
	8'h75: num[23:16] = 8'hd3;
	8'h76: num[23:16] = 8'h27;
	8'h77: num[23:16] = 8'h52;
	8'h78: num[23:16] = 8'h4c;
	8'h79: num[23:16] = 8'h36;
	8'h7a: num[23:16] = 8'h02;
	8'h7b: num[23:16] = 8'he7;
	8'h7c: num[23:16] = 8'ha0;
	8'h7d: num[23:16] = 8'hc4;
	8'h7e: num[23:16] = 8'hc8;
	8'h7f: num[23:16] = 8'h9e;
	8'h80: num[23:16] = 8'hea;
	8'h81: num[23:16] = 8'hbf;
	8'h82: num[23:16] = 8'h8a;
	8'h83: num[23:16] = 8'hd2;
	8'h84: num[23:16] = 8'h40;
	8'h85: num[23:16] = 8'hc7;
	8'h86: num[23:16] = 8'h38;
	8'h87: num[23:16] = 8'hb5;
	8'h88: num[23:16] = 8'ha3;
	8'h89: num[23:16] = 8'hf7;
	8'h8a: num[23:16] = 8'hf2;
	8'h8b: num[23:16] = 8'hce;
	8'h8c: num[23:16] = 8'hf9;
	8'h8d: num[23:16] = 8'h61;
	8'h8e: num[23:16] = 8'h15;
	8'h8f: num[23:16] = 8'ha1;
	8'h90: num[23:16] = 8'he0;
	8'h91: num[23:16] = 8'hae;
	8'h92: num[23:16] = 8'h5d;
	8'h93: num[23:16] = 8'ha4;
	8'h94: num[23:16] = 8'h9b;
	8'h95: num[23:16] = 8'h34;
	8'h96: num[23:16] = 8'h1a;
	8'h97: num[23:16] = 8'h55;
	8'h98: num[23:16] = 8'had;
	8'h99: num[23:16] = 8'h93;
	8'h9a: num[23:16] = 8'h32;
	8'h9b: num[23:16] = 8'h30;
	8'h9c: num[23:16] = 8'hf5;
	8'h9d: num[23:16] = 8'h8c;
	8'h9e: num[23:16] = 8'hb1;
	8'h9f: num[23:16] = 8'he3;
	8'ha0: num[23:16] = 8'h1d;
	8'ha1: num[23:16] = 8'hf6;
	8'ha2: num[23:16] = 8'he2;
	8'ha3: num[23:16] = 8'h2e;
	8'ha4: num[23:16] = 8'h82;
	8'ha5: num[23:16] = 8'h66;
	8'ha6: num[23:16] = 8'hca;
	8'ha7: num[23:16] = 8'h60;
	8'ha8: num[23:16] = 8'hc0;
	8'ha9: num[23:16] = 8'h29;
	8'haa: num[23:16] = 8'h23;
	8'hab: num[23:16] = 8'hab;
	8'hac: num[23:16] = 8'h0d;
	8'had: num[23:16] = 8'h53;
	8'hae: num[23:16] = 8'h4e;
	8'haf: num[23:16] = 8'h6f;
	8'hb0: num[23:16] = 8'hd5;
	8'hb1: num[23:16] = 8'hdb;
	8'hb2: num[23:16] = 8'h37;
	8'hb3: num[23:16] = 8'h45;
	8'hb4: num[23:16] = 8'hde;
	8'hb5: num[23:16] = 8'hfd;
	8'hb6: num[23:16] = 8'h8e;
	8'hb7: num[23:16] = 8'h2f;
	8'hb8: num[23:16] = 8'h03;
	8'hb9: num[23:16] = 8'hff;
	8'hba: num[23:16] = 8'h6a;
	8'hbb: num[23:16] = 8'h72;
	8'hbc: num[23:16] = 8'h6d;
	8'hbd: num[23:16] = 8'h6c;
	8'hbe: num[23:16] = 8'h5b;
	8'hbf: num[23:16] = 8'h51;
	8'hc0: num[23:16] = 8'h8d;
	8'hc1: num[23:16] = 8'h1b;
	8'hc2: num[23:16] = 8'haf;
	8'hc3: num[23:16] = 8'h92;
	8'hc4: num[23:16] = 8'hbb;
	8'hc5: num[23:16] = 8'hdd;
	8'hc6: num[23:16] = 8'hbc;
	8'hc7: num[23:16] = 8'h7f;
	8'hc8: num[23:16] = 8'h11;
	8'hc9: num[23:16] = 8'hd9;
	8'hca: num[23:16] = 8'h5c;
	8'hcb: num[23:16] = 8'h41;
	8'hcc: num[23:16] = 8'h1f;
	8'hcd: num[23:16] = 8'h10;
	8'hce: num[23:16] = 8'h5a;
	8'hcf: num[23:16] = 8'hd8;
	8'hd0: num[23:16] = 8'h0a;
	8'hd1: num[23:16] = 8'hc1;
	8'hd2: num[23:16] = 8'h31;
	8'hd3: num[23:16] = 8'h88;
	8'hd4: num[23:16] = 8'ha5;
	8'hd5: num[23:16] = 8'hcd;
	8'hd6: num[23:16] = 8'h7b;
	8'hd7: num[23:16] = 8'hbd;
	8'hd8: num[23:16] = 8'h2d;
	8'hd9: num[23:16] = 8'h74;
	8'hda: num[23:16] = 8'hd0;
	8'hdb: num[23:16] = 8'h12;
	8'hdc: num[23:16] = 8'hb8;
	8'hdd: num[23:16] = 8'he5;
	8'hde: num[23:16] = 8'hb4;
	8'hdf: num[23:16] = 8'hb0;
	8'he0: num[23:16] = 8'h89;
	8'he1: num[23:16] = 8'h69;
	8'he2: num[23:16] = 8'h97;
	8'he3: num[23:16] = 8'h4a;
	8'he4: num[23:16] = 8'h0c;
	8'he5: num[23:16] = 8'h96;
	8'he6: num[23:16] = 8'h77;
	8'he7: num[23:16] = 8'h7e;
	8'he8: num[23:16] = 8'h65;
	8'he9: num[23:16] = 8'hb9;
	8'hea: num[23:16] = 8'hf1;
	8'heb: num[23:16] = 8'h09;
	8'hec: num[23:16] = 8'hc5;
	8'hed: num[23:16] = 8'h6e;
	8'hee: num[23:16] = 8'hc6;
	8'hef: num[23:16] = 8'h84;
	8'hf0: num[23:16] = 8'h18;
	8'hf1: num[23:16] = 8'hf0;
	8'hf2: num[23:16] = 8'h7d;
	8'hf3: num[23:16] = 8'hec;
	8'hf4: num[23:16] = 8'h3a;
	8'hf5: num[23:16] = 8'hdc;
	8'hf6: num[23:16] = 8'h4d;
	8'hf7: num[23:16] = 8'h20;
	8'hf8: num[23:16] = 8'h79;
	8'hf9: num[23:16] = 8'hee;
	8'hfa: num[23:16] = 8'h5f;
	8'hfb: num[23:16] = 8'h3e;
	8'hfc: num[23:16] = 8'hd7;
	8'hfd: num[23:16] = 8'hcb;
	8'hfe: num[23:16] = 8'h39;
	8'hff: num[23:16] = 8'h48;
	default: num[23:16] = 8'h00;
	endcase
	case(num[31:24])
	8'h00: num[31:24] = 8'hd6;
	8'h01: num[31:24] = 8'h90;
	8'h02: num[31:24] = 8'he9;
	8'h03: num[31:24] = 8'hfe;
	8'h04: num[31:24] = 8'hcc;
	8'h05: num[31:24] = 8'he1;
	8'h06: num[31:24] = 8'h3d;
	8'h07: num[31:24] = 8'hb7;
	8'h08: num[31:24] = 8'h16;
	8'h09: num[31:24] = 8'hb6;
	8'h0a: num[31:24] = 8'h14;
	8'h0b: num[31:24] = 8'hc2;
	8'h0c: num[31:24] = 8'h28;
	8'h0d: num[31:24] = 8'hfb;
	8'h0e: num[31:24] = 8'h2c;
	8'h0f: num[31:24] = 8'h05;
	8'h10: num[31:24] = 8'h2b;
	8'h11: num[31:24] = 8'h67;
	8'h12: num[31:24] = 8'h9a;
	8'h13: num[31:24] = 8'h76;
	8'h14: num[31:24] = 8'h2a;
	8'h15: num[31:24] = 8'hbe;
	8'h16: num[31:24] = 8'h04;
	8'h17: num[31:24] = 8'hc3;
	8'h18: num[31:24] = 8'haa;
	8'h19: num[31:24] = 8'h44;
	8'h1a: num[31:24] = 8'h13;
	8'h1b: num[31:24] = 8'h26;
	8'h1c: num[31:24] = 8'h49;
	8'h1d: num[31:24] = 8'h86;
	8'h1e: num[31:24] = 8'h06;
	8'h1f: num[31:24] = 8'h99;
	8'h20: num[31:24] = 8'h9c;
	8'h21: num[31:24] = 8'h42;
	8'h22: num[31:24] = 8'h50;
	8'h23: num[31:24] = 8'hf4;
	8'h24: num[31:24] = 8'h91;
	8'h25: num[31:24] = 8'hef;
	8'h26: num[31:24] = 8'h98;
	8'h27: num[31:24] = 8'h7a;
	8'h28: num[31:24] = 8'h33;
	8'h29: num[31:24] = 8'h54;
	8'h2a: num[31:24] = 8'h0b;
	8'h2b: num[31:24] = 8'h43;
	8'h2c: num[31:24] = 8'hed;
	8'h2d: num[31:24] = 8'hcf;
	8'h2e: num[31:24] = 8'hac;
	8'h2f: num[31:24] = 8'h62;
	8'h30: num[31:24] = 8'he4;
	8'h31: num[31:24] = 8'hb3;
	8'h32: num[31:24] = 8'h1c;
	8'h33: num[31:24] = 8'ha9;
	8'h34: num[31:24] = 8'hc9;
	8'h35: num[31:24] = 8'h08;
	8'h36: num[31:24] = 8'he8;
	8'h37: num[31:24] = 8'h95;
	8'h38: num[31:24] = 8'h80;
	8'h39: num[31:24] = 8'hdf;
	8'h3a: num[31:24] = 8'h94;
	8'h3b: num[31:24] = 8'hfa;
	8'h3c: num[31:24] = 8'h75;
	8'h3d: num[31:24] = 8'h8f;
	8'h3e: num[31:24] = 8'h3f;
	8'h3f: num[31:24] = 8'ha6;
	8'h40: num[31:24] = 8'h47;
	8'h41: num[31:24] = 8'h07;
	8'h42: num[31:24] = 8'ha7;
	8'h43: num[31:24] = 8'hfc;
	8'h44: num[31:24] = 8'hf3;
	8'h45: num[31:24] = 8'h73;
	8'h46: num[31:24] = 8'h17;
	8'h47: num[31:24] = 8'hba;
	8'h48: num[31:24] = 8'h83;
	8'h49: num[31:24] = 8'h59;
	8'h4a: num[31:24] = 8'h3c;
	8'h4b: num[31:24] = 8'h19;
	8'h4c: num[31:24] = 8'he6;
	8'h4d: num[31:24] = 8'h85;
	8'h4e: num[31:24] = 8'h4f;
	8'h4f: num[31:24] = 8'ha8;
	8'h50: num[31:24] = 8'h68;
	8'h51: num[31:24] = 8'h6b;
	8'h52: num[31:24] = 8'h81;
	8'h53: num[31:24] = 8'hb2;
	8'h54: num[31:24] = 8'h71;
	8'h55: num[31:24] = 8'h64;
	8'h56: num[31:24] = 8'hda;
	8'h57: num[31:24] = 8'h8b;
	8'h58: num[31:24] = 8'hf8;
	8'h59: num[31:24] = 8'heb;
	8'h5a: num[31:24] = 8'h0f;
	8'h5b: num[31:24] = 8'h4b;
	8'h5c: num[31:24] = 8'h70;
	8'h5d: num[31:24] = 8'h56;
	8'h5e: num[31:24] = 8'h9d;
	8'h5f: num[31:24] = 8'h35;
	8'h60: num[31:24] = 8'h1e;
	8'h61: num[31:24] = 8'h24;
	8'h62: num[31:24] = 8'h0e;
	8'h63: num[31:24] = 8'h5e;
	8'h64: num[31:24] = 8'h63;
	8'h65: num[31:24] = 8'h58;
	8'h66: num[31:24] = 8'hd1;
	8'h67: num[31:24] = 8'ha2;
	8'h68: num[31:24] = 8'h25;
	8'h69: num[31:24] = 8'h22;
	8'h6a: num[31:24] = 8'h7c;
	8'h6b: num[31:24] = 8'h3b;
	8'h6c: num[31:24] = 8'h01;
	8'h6d: num[31:24] = 8'h21;
	8'h6e: num[31:24] = 8'h78;
	8'h6f: num[31:24] = 8'h87;
	8'h70: num[31:24] = 8'hd4;
	8'h71: num[31:24] = 8'h00;
	8'h72: num[31:24] = 8'h46;
	8'h73: num[31:24] = 8'h57;
	8'h74: num[31:24] = 8'h9f;
	8'h75: num[31:24] = 8'hd3;
	8'h76: num[31:24] = 8'h27;
	8'h77: num[31:24] = 8'h52;
	8'h78: num[31:24] = 8'h4c;
	8'h79: num[31:24] = 8'h36;
	8'h7a: num[31:24] = 8'h02;
	8'h7b: num[31:24] = 8'he7;
	8'h7c: num[31:24] = 8'ha0;
	8'h7d: num[31:24] = 8'hc4;
	8'h7e: num[31:24] = 8'hc8;
	8'h7f: num[31:24] = 8'h9e;
	8'h80: num[31:24] = 8'hea;
	8'h81: num[31:24] = 8'hbf;
	8'h82: num[31:24] = 8'h8a;
	8'h83: num[31:24] = 8'hd2;
	8'h84: num[31:24] = 8'h40;
	8'h85: num[31:24] = 8'hc7;
	8'h86: num[31:24] = 8'h38;
	8'h87: num[31:24] = 8'hb5;
	8'h88: num[31:24] = 8'ha3;
	8'h89: num[31:24] = 8'hf7;
	8'h8a: num[31:24] = 8'hf2;
	8'h8b: num[31:24] = 8'hce;
	8'h8c: num[31:24] = 8'hf9;
	8'h8d: num[31:24] = 8'h61;
	8'h8e: num[31:24] = 8'h15;
	8'h8f: num[31:24] = 8'ha1;
	8'h90: num[31:24] = 8'he0;
	8'h91: num[31:24] = 8'hae;
	8'h92: num[31:24] = 8'h5d;
	8'h93: num[31:24] = 8'ha4;
	8'h94: num[31:24] = 8'h9b;
	8'h95: num[31:24] = 8'h34;
	8'h96: num[31:24] = 8'h1a;
	8'h97: num[31:24] = 8'h55;
	8'h98: num[31:24] = 8'had;
	8'h99: num[31:24] = 8'h93;
	8'h9a: num[31:24] = 8'h32;
	8'h9b: num[31:24] = 8'h30;
	8'h9c: num[31:24] = 8'hf5;
	8'h9d: num[31:24] = 8'h8c;
	8'h9e: num[31:24] = 8'hb1;
	8'h9f: num[31:24] = 8'he3;
	8'ha0: num[31:24] = 8'h1d;
	8'ha1: num[31:24] = 8'hf6;
	8'ha2: num[31:24] = 8'he2;
	8'ha3: num[31:24] = 8'h2e;
	8'ha4: num[31:24] = 8'h82;
	8'ha5: num[31:24] = 8'h66;
	8'ha6: num[31:24] = 8'hca;
	8'ha7: num[31:24] = 8'h60;
	8'ha8: num[31:24] = 8'hc0;
	8'ha9: num[31:24] = 8'h29;
	8'haa: num[31:24] = 8'h23;
	8'hab: num[31:24] = 8'hab;
	8'hac: num[31:24] = 8'h0d;
	8'had: num[31:24] = 8'h53;
	8'hae: num[31:24] = 8'h4e;
	8'haf: num[31:24] = 8'h6f;
	8'hb0: num[31:24] = 8'hd5;
	8'hb1: num[31:24] = 8'hdb;
	8'hb2: num[31:24] = 8'h37;
	8'hb3: num[31:24] = 8'h45;
	8'hb4: num[31:24] = 8'hde;
	8'hb5: num[31:24] = 8'hfd;
	8'hb6: num[31:24] = 8'h8e;
	8'hb7: num[31:24] = 8'h2f;
	8'hb8: num[31:24] = 8'h03;
	8'hb9: num[31:24] = 8'hff;
	8'hba: num[31:24] = 8'h6a;
	8'hbb: num[31:24] = 8'h72;
	8'hbc: num[31:24] = 8'h6d;
	8'hbd: num[31:24] = 8'h6c;
	8'hbe: num[31:24] = 8'h5b;
	8'hbf: num[31:24] = 8'h51;
	8'hc0: num[31:24] = 8'h8d;
	8'hc1: num[31:24] = 8'h1b;
	8'hc2: num[31:24] = 8'haf;
	8'hc3: num[31:24] = 8'h92;
	8'hc4: num[31:24] = 8'hbb;
	8'hc5: num[31:24] = 8'hdd;
	8'hc6: num[31:24] = 8'hbc;
	8'hc7: num[31:24] = 8'h7f;
	8'hc8: num[31:24] = 8'h11;
	8'hc9: num[31:24] = 8'hd9;
	8'hca: num[31:24] = 8'h5c;
	8'hcb: num[31:24] = 8'h41;
	8'hcc: num[31:24] = 8'h1f;
	8'hcd: num[31:24] = 8'h10;
	8'hce: num[31:24] = 8'h5a;
	8'hcf: num[31:24] = 8'hd8;
	8'hd0: num[31:24] = 8'h0a;
	8'hd1: num[31:24] = 8'hc1;
	8'hd2: num[31:24] = 8'h31;
	8'hd3: num[31:24] = 8'h88;
	8'hd4: num[31:24] = 8'ha5;
	8'hd5: num[31:24] = 8'hcd;
	8'hd6: num[31:24] = 8'h7b;
	8'hd7: num[31:24] = 8'hbd;
	8'hd8: num[31:24] = 8'h2d;
	8'hd9: num[31:24] = 8'h74;
	8'hda: num[31:24] = 8'hd0;
	8'hdb: num[31:24] = 8'h12;
	8'hdc: num[31:24] = 8'hb8;
	8'hdd: num[31:24] = 8'he5;
	8'hde: num[31:24] = 8'hb4;
	8'hdf: num[31:24] = 8'hb0;
	8'he0: num[31:24] = 8'h89;
	8'he1: num[31:24] = 8'h69;
	8'he2: num[31:24] = 8'h97;
	8'he3: num[31:24] = 8'h4a;
	8'he4: num[31:24] = 8'h0c;
	8'he5: num[31:24] = 8'h96;
	8'he6: num[31:24] = 8'h77;
	8'he7: num[31:24] = 8'h7e;
	8'he8: num[31:24] = 8'h65;
	8'he9: num[31:24] = 8'hb9;
	8'hea: num[31:24] = 8'hf1;
	8'heb: num[31:24] = 8'h09;
	8'hec: num[31:24] = 8'hc5;
	8'hed: num[31:24] = 8'h6e;
	8'hee: num[31:24] = 8'hc6;
	8'hef: num[31:24] = 8'h84;
	8'hf0: num[31:24] = 8'h18;
	8'hf1: num[31:24] = 8'hf0;
	8'hf2: num[31:24] = 8'h7d;
	8'hf3: num[31:24] = 8'hec;
	8'hf4: num[31:24] = 8'h3a;
	8'hf5: num[31:24] = 8'hdc;
	8'hf6: num[31:24] = 8'h4d;
	8'hf7: num[31:24] = 8'h20;
	8'hf8: num[31:24] = 8'h79;
	8'hf9: num[31:24] = 8'hee;
	8'hfa: num[31:24] = 8'h5f;
	8'hfb: num[31:24] = 8'h3e;
	8'hfc: num[31:24] = 8'hd7;
	8'hfd: num[31:24] = 8'hcb;
	8'hfe: num[31:24] = 8'h39;
	8'hff: num[31:24] = 8'h48;
	default: num[31:24] = 8'h00;
	endcase
	text[i+4] = text[i] ^ num ^ {num[29:0], num[31:30]} ^ {num[21:0], num[31:22]} ^ {num[13:0], num[31:14]} ^ {num[7:0],num[31:8]};
	
	cipher = {text[35], text[34], text[33], text[32]};
    end
    
    end
    
    
    
    
endmodule